magic
tech s8seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
rect 410 2294 470 51210
tri 410 2269 470 2294 nw
<< end >>
