# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_io__top_gpiov2
  CLASS PAD ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 80 BY 200 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 53.125000 1.270000 56.105000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 53.125000 80.000000 56.105000 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    ANTENNAPARTIALMETALSIDEAREA  119.1680 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000000 48.365000 1.270000 51.345000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 48.365000 80.000000 51.345000 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430000 0.000000 62.690000 1.915000 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865000  0.000000 46.195000 36.665000 ;
        RECT 45.865000 36.665000 46.195000 36.735000 ;
        RECT 45.865000 36.735000 46.265000 36.805000 ;
        RECT 45.965000 36.805000 46.335000 36.905000 ;
        RECT 46.065000 36.905000 46.435000 37.005000 ;
        RECT 46.070000 37.005000 46.535000 37.010000 ;
        RECT 46.220000 37.010000 48.225000 37.160000 ;
        RECT 46.370000 37.160000 48.075000 37.310000 ;
        RECT 46.400000 37.310000 48.045000 37.340000 ;
        RECT 47.910000 37.005000 48.375000 37.010000 ;
        RECT 47.960000 35.870000 48.740000 36.190000 ;
        RECT 47.975000 36.940000 48.380000 37.005000 ;
        RECT 48.040000 36.875000 48.445000 36.940000 ;
        RECT 48.070000 36.190000 48.630000 36.300000 ;
        RECT 48.110000 36.805000 48.510000 36.875000 ;
        RECT 48.180000 36.300000 48.520000 36.410000 ;
        RECT 48.180000 36.410000 48.515000 36.415000 ;
        RECT 48.180000 36.415000 48.510000 36.420000 ;
        RECT 48.180000 36.420000 48.510000 36.735000 ;
        RECT 48.180000 36.735000 48.510000 36.805000 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.080000 57.360000 24.590000 57.430000 ;
        RECT 23.080000 57.430000 24.520000 57.500000 ;
        RECT 23.080000 57.500000 24.450000 57.570000 ;
        RECT 23.080000 57.570000 24.380000 57.640000 ;
        RECT 24.285000 57.345000 24.660000 57.360000 ;
        RECT 24.355000 57.275000 24.675000 57.345000 ;
        RECT 24.425000 57.205000 24.745000 57.275000 ;
        RECT 24.495000 57.135000 24.815000 57.205000 ;
        RECT 24.565000 57.065000 24.885000 57.135000 ;
        RECT 24.620000 57.010000 24.955000 57.065000 ;
        RECT 24.675000 53.255000 25.010000 53.310000 ;
        RECT 24.675000 53.310000 24.955000 53.365000 ;
        RECT 24.675000 53.365000 24.955000 56.955000 ;
        RECT 24.675000 56.955000 24.955000 57.010000 ;
        RECT 24.740000 53.190000 25.065000 53.255000 ;
        RECT 24.810000 53.120000 25.130000 53.190000 ;
        RECT 24.880000 53.050000 25.200000 53.120000 ;
        RECT 24.950000 52.980000 25.270000 53.050000 ;
        RECT 25.020000 52.910000 25.340000 52.980000 ;
        RECT 25.090000 52.840000 25.410000 52.910000 ;
        RECT 25.160000 52.770000 25.480000 52.840000 ;
        RECT 25.230000 52.700000 25.550000 52.770000 ;
        RECT 25.300000 52.630000 25.620000 52.700000 ;
        RECT 25.370000 52.560000 25.690000 52.630000 ;
        RECT 25.440000 52.490000 25.760000 52.560000 ;
        RECT 25.510000 52.420000 25.830000 52.490000 ;
        RECT 25.580000 52.350000 25.900000 52.420000 ;
        RECT 25.650000 52.280000 25.970000 52.350000 ;
        RECT 25.720000 52.210000 26.040000 52.280000 ;
        RECT 25.790000 52.140000 29.735000 52.210000 ;
        RECT 25.860000 52.070000 29.805000 52.140000 ;
        RECT 25.930000 52.000000 29.875000 52.070000 ;
        RECT 26.000000 51.930000 29.945000 52.000000 ;
        RECT 29.645000 51.910000 30.015000 51.930000 ;
        RECT 29.715000 51.840000 30.035000 51.910000 ;
        RECT 29.785000 51.770000 30.105000 51.840000 ;
        RECT 29.855000 51.700000 30.175000 51.770000 ;
        RECT 29.925000 51.630000 30.245000 51.700000 ;
        RECT 29.995000 51.560000 30.315000 51.630000 ;
        RECT 30.060000 51.495000 30.385000 51.560000 ;
        RECT 30.125000 17.630000 30.440000 17.685000 ;
        RECT 30.125000 17.685000 30.385000 17.740000 ;
        RECT 30.125000 17.740000 30.385000 36.345000 ;
        RECT 30.125000 36.345000 30.385000 36.400000 ;
        RECT 30.125000 36.400000 30.440000 36.455000 ;
        RECT 30.125000 38.010000 30.440000 38.065000 ;
        RECT 30.125000 38.065000 30.385000 38.120000 ;
        RECT 30.125000 38.120000 30.385000 51.430000 ;
        RECT 30.125000 51.430000 30.385000 51.495000 ;
        RECT 30.140000 37.995000 30.495000 38.010000 ;
        RECT 30.180000 17.575000 30.495000 17.630000 ;
        RECT 30.195000 36.455000 30.495000 36.525000 ;
        RECT 30.210000 37.925000 30.510000 37.995000 ;
        RECT 30.250000 17.505000 30.550000 17.575000 ;
        RECT 30.265000 36.525000 30.565000 36.595000 ;
        RECT 30.280000 36.595000 30.635000 36.610000 ;
        RECT 30.280000 37.855000 30.580000 37.925000 ;
        RECT 30.320000 17.435000 30.620000 17.505000 ;
        RECT 30.335000 36.610000 30.650000 36.665000 ;
        RECT 30.335000 37.800000 30.650000 37.855000 ;
        RECT 30.390000 17.365000 30.690000 17.435000 ;
        RECT 30.390000 36.665000 30.650000 36.720000 ;
        RECT 30.390000 36.720000 30.650000 37.745000 ;
        RECT 30.390000 37.745000 30.650000 37.800000 ;
        RECT 30.460000 17.295000 30.760000 17.365000 ;
        RECT 30.530000 17.225000 30.830000 17.295000 ;
        RECT 30.600000 17.155000 30.900000 17.225000 ;
        RECT 30.670000 17.085000 30.970000 17.155000 ;
        RECT 30.740000 17.015000 31.040000 17.085000 ;
        RECT 30.750000  0.000000 31.010000  2.155000 ;
        RECT 30.750000  2.155000 31.010000  2.210000 ;
        RECT 30.750000  2.210000 31.065000  2.265000 ;
        RECT 30.810000 16.945000 31.110000 17.015000 ;
        RECT 30.820000  2.265000 31.120000  2.335000 ;
        RECT 30.880000 16.875000 31.180000 16.945000 ;
        RECT 30.890000  2.335000 31.190000  2.405000 ;
        RECT 30.950000 16.805000 31.250000 16.875000 ;
        RECT 30.960000  2.405000 31.260000  2.475000 ;
        RECT 31.020000 16.735000 31.320000 16.805000 ;
        RECT 31.030000  2.475000 31.330000  2.545000 ;
        RECT 31.090000 16.665000 31.390000 16.735000 ;
        RECT 31.100000  2.545000 31.400000  2.615000 ;
        RECT 31.160000 16.595000 31.460000 16.665000 ;
        RECT 31.170000  2.615000 31.470000  2.685000 ;
        RECT 31.195000  2.685000 31.540000  2.710000 ;
        RECT 31.230000 16.525000 31.530000 16.595000 ;
        RECT 31.250000  2.710000 31.565000  2.765000 ;
        RECT 31.300000 16.455000 31.600000 16.525000 ;
        RECT 31.305000  2.765000 31.565000  2.820000 ;
        RECT 31.305000  2.820000 31.565000  4.335000 ;
        RECT 31.305000  4.335000 31.565000  4.390000 ;
        RECT 31.305000  4.390000 31.620000  4.445000 ;
        RECT 31.370000 16.385000 31.670000 16.455000 ;
        RECT 31.375000  4.445000 31.675000  4.515000 ;
        RECT 31.440000 16.315000 31.740000 16.385000 ;
        RECT 31.445000  4.515000 31.745000  4.585000 ;
        RECT 31.510000 16.245000 31.810000 16.315000 ;
        RECT 31.515000  4.585000 31.815000  4.655000 ;
        RECT 31.580000  4.655000 31.885000  4.720000 ;
        RECT 31.580000 16.175000 31.880000 16.245000 ;
        RECT 31.635000  4.720000 31.950000  4.775000 ;
        RECT 31.635000 16.120000 31.950000 16.175000 ;
        RECT 31.690000  4.775000 31.950000  4.830000 ;
        RECT 31.690000  4.830000 31.950000 16.065000 ;
        RECT 31.690000 16.065000 31.950000 16.120000 ;
    END
  END ANALOG_SEL
  PIN DM[0]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.590000 0.545000 50.360000 0.825000 ;
        RECT 49.625000 0.510000 50.325000 0.545000 ;
        RECT 49.695000 0.440000 50.255000 0.510000 ;
        RECT 49.765000 0.370000 50.185000 0.440000 ;
        RECT 49.835000 0.300000 50.115000 0.370000 ;
        RECT 49.845000 0.290000 50.115000 0.300000 ;
        RECT 49.855000 0.000000 50.115000 0.280000 ;
        RECT 49.855000 0.280000 50.115000 0.290000 ;
    END
  END DM[0]
  PIN DM[1]
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.540000 1.195000 67.360000 1.475000 ;
        RECT 66.595000 1.140000 67.305000 1.195000 ;
        RECT 66.665000 1.070000 67.235000 1.140000 ;
        RECT 66.735000 1.000000 67.165000 1.070000 ;
        RECT 66.805000 0.930000 67.095000 1.000000 ;
        RECT 66.820000 0.915000 67.095000 0.930000 ;
        RECT 66.835000 0.000000 67.095000 0.900000 ;
        RECT 66.835000 0.900000 67.095000 0.915000 ;
    END
  END DM[1]
  PIN DM[2]
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490000 0.000000 28.750000 3.960000 ;
        RECT 28.490000 3.960000 28.750000 4.015000 ;
        RECT 28.490000 4.015000 28.805000 4.070000 ;
        RECT 28.560000 4.070000 28.860000 4.140000 ;
        RECT 28.630000 4.140000 28.930000 4.210000 ;
        RECT 28.700000 4.210000 29.000000 4.280000 ;
        RECT 28.770000 4.280000 29.070000 4.350000 ;
        RECT 28.840000 4.350000 29.140000 4.420000 ;
        RECT 28.910000 4.420000 29.210000 4.490000 ;
        RECT 28.980000 4.490000 29.280000 4.560000 ;
        RECT 29.050000 4.560000 29.350000 4.630000 ;
        RECT 29.100000 4.630000 29.420000 4.680000 ;
        RECT 29.155000 4.680000 29.470000 4.735000 ;
        RECT 29.210000 4.735000 29.470000 4.790000 ;
        RECT 29.210000 4.790000 29.470000 6.780000 ;
    END
  END DM[2]
  PIN ENABLE_H
    ANTENNAGATEAREA  4.860000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.135000 2.225000 35.450000 2.280000 ;
        RECT 35.135000 2.280000 35.395000 2.335000 ;
        RECT 35.135000 2.335000 35.395000 3.885000 ;
        RECT 35.140000 2.220000 35.505000 2.225000 ;
        RECT 35.210000 2.150000 35.510000 2.220000 ;
        RECT 35.280000 2.080000 35.580000 2.150000 ;
        RECT 35.350000 2.010000 35.650000 2.080000 ;
        RECT 35.405000 1.955000 35.720000 2.010000 ;
        RECT 35.460000 0.000000 35.720000 1.900000 ;
        RECT 35.460000 1.900000 35.720000 1.955000 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390000 0.000000 38.650000 3.715000 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    ANTENNAGATEAREA  3.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.315000 56.460000  7.630000 56.515000 ;
        RECT  7.315000 56.515000  7.575000 56.570000 ;
        RECT  7.315000 56.570000  7.575000 73.615000 ;
        RECT  7.315000 73.615000  7.575000 73.670000 ;
        RECT  7.315000 73.670000  7.630000 73.725000 ;
        RECT  7.375000 56.400000  7.685000 56.460000 ;
        RECT  7.385000 73.725000  7.685000 73.795000 ;
        RECT  7.445000 56.330000  7.745000 56.400000 ;
        RECT  7.455000 73.795000  7.755000 73.865000 ;
        RECT  7.515000 56.260000  7.815000 56.330000 ;
        RECT  7.525000 73.865000  7.825000 73.935000 ;
        RECT  7.585000 56.190000  7.885000 56.260000 ;
        RECT  7.595000 73.935000  7.895000 74.005000 ;
        RECT  7.655000 56.120000  7.955000 56.190000 ;
        RECT  7.665000 74.005000  7.965000 74.075000 ;
        RECT  7.695000 74.075000  8.035000 74.105000 ;
        RECT  7.725000 56.050000  8.025000 56.120000 ;
        RECT  7.750000 74.105000  8.065000 74.160000 ;
        RECT  7.795000 55.980000  8.095000 56.050000 ;
        RECT  7.805000 74.160000  8.065000 74.215000 ;
        RECT  7.805000 74.215000  8.065000 74.680000 ;
        RECT  7.805000 74.680000  8.065000 74.735000 ;
        RECT  7.805000 74.735000  8.120000 74.790000 ;
        RECT  7.865000 55.910000  8.165000 55.980000 ;
        RECT  7.875000 74.790000  8.175000 74.860000 ;
        RECT  7.920000 55.855000  8.235000 55.910000 ;
        RECT  7.920000 77.285000  8.560000 77.545000 ;
        RECT  7.945000 74.860000  8.245000 74.930000 ;
        RECT  7.975000 53.960000  8.290000 54.015000 ;
        RECT  7.975000 54.015000  8.235000 54.070000 ;
        RECT  7.975000 54.070000  8.235000 55.800000 ;
        RECT  7.975000 55.800000  8.235000 55.855000 ;
        RECT  8.015000 74.930000  8.315000 75.000000 ;
        RECT  8.030000 53.905000  8.345000 53.960000 ;
        RECT  8.085000 53.850000  8.400000 53.905000 ;
        RECT  8.085000 75.000000  8.385000 75.070000 ;
        RECT  8.085000 77.240000  8.515000 77.285000 ;
        RECT  8.100000 75.070000  8.455000 75.085000 ;
        RECT  8.130000 77.195000  8.470000 77.240000 ;
        RECT  8.140000 53.795000  8.455000 53.850000 ;
        RECT  8.155000 75.085000  8.470000 75.140000 ;
        RECT  8.170000 77.155000  8.470000 77.195000 ;
        RECT  8.195000 44.075000  8.510000 44.130000 ;
        RECT  8.195000 44.130000  8.455000 44.185000 ;
        RECT  8.195000 44.185000  8.455000 53.740000 ;
        RECT  8.195000 53.740000  8.455000 53.795000 ;
        RECT  8.210000 44.060000  8.565000 44.075000 ;
        RECT  8.210000 75.140000  8.470000 75.195000 ;
        RECT  8.210000 75.195000  8.470000 77.115000 ;
        RECT  8.210000 77.115000  8.470000 77.155000 ;
        RECT  8.280000 43.990000  8.580000 44.060000 ;
        RECT  8.350000 43.920000  8.650000 43.990000 ;
        RECT  8.420000 43.850000  8.720000 43.920000 ;
        RECT  8.490000 43.780000  8.790000 43.850000 ;
        RECT  8.560000 43.710000  8.860000 43.780000 ;
        RECT  8.630000 43.640000  8.930000 43.710000 ;
        RECT  8.700000 43.570000  9.000000 43.640000 ;
        RECT  8.770000 43.500000  9.070000 43.570000 ;
        RECT  8.840000 43.430000  9.140000 43.500000 ;
        RECT  8.910000 43.360000  9.210000 43.430000 ;
        RECT  8.980000 43.290000  9.280000 43.360000 ;
        RECT  9.050000 43.220000  9.350000 43.290000 ;
        RECT  9.120000 43.150000  9.420000 43.220000 ;
        RECT  9.190000 43.080000  9.490000 43.150000 ;
        RECT  9.260000 43.010000  9.560000 43.080000 ;
        RECT  9.330000 42.940000  9.630000 43.010000 ;
        RECT  9.400000 42.870000  9.700000 42.940000 ;
        RECT  9.470000 42.800000  9.770000 42.870000 ;
        RECT  9.540000 42.730000  9.840000 42.800000 ;
        RECT  9.610000 42.660000  9.910000 42.730000 ;
        RECT  9.680000 42.590000  9.980000 42.660000 ;
        RECT  9.750000 42.520000 10.050000 42.590000 ;
        RECT  9.820000 42.450000 10.120000 42.520000 ;
        RECT  9.890000 42.380000 10.190000 42.450000 ;
        RECT  9.960000 42.310000 10.260000 42.380000 ;
        RECT 10.030000 42.240000 10.330000 42.310000 ;
        RECT 10.100000 42.170000 10.400000 42.240000 ;
        RECT 10.170000 42.100000 10.470000 42.170000 ;
        RECT 10.240000 42.030000 10.540000 42.100000 ;
        RECT 10.310000 41.960000 10.610000 42.030000 ;
        RECT 10.380000 41.890000 10.680000 41.960000 ;
        RECT 10.450000 41.820000 10.750000 41.890000 ;
        RECT 10.520000 41.750000 10.820000 41.820000 ;
        RECT 10.590000 41.680000 10.890000 41.750000 ;
        RECT 10.660000 41.610000 10.960000 41.680000 ;
        RECT 10.730000 41.540000 11.030000 41.610000 ;
        RECT 10.800000 41.470000 11.100000 41.540000 ;
        RECT 10.870000 41.400000 11.170000 41.470000 ;
        RECT 10.940000 41.330000 11.240000 41.400000 ;
        RECT 11.010000 41.260000 11.310000 41.330000 ;
        RECT 11.080000 41.190000 11.380000 41.260000 ;
        RECT 11.150000 41.120000 11.450000 41.190000 ;
        RECT 11.220000 41.050000 11.520000 41.120000 ;
        RECT 11.290000 40.980000 11.590000 41.050000 ;
        RECT 11.360000 40.910000 11.660000 40.980000 ;
        RECT 11.430000 40.840000 11.730000 40.910000 ;
        RECT 11.500000 40.770000 11.800000 40.840000 ;
        RECT 11.570000 40.700000 11.870000 40.770000 ;
        RECT 11.640000 40.630000 11.940000 40.700000 ;
        RECT 11.710000 40.560000 12.010000 40.630000 ;
        RECT 11.780000 40.490000 12.080000 40.560000 ;
        RECT 11.850000 40.420000 12.150000 40.490000 ;
        RECT 11.920000 40.350000 12.220000 40.420000 ;
        RECT 11.990000 40.280000 12.290000 40.350000 ;
        RECT 12.060000 40.210000 12.360000 40.280000 ;
        RECT 12.130000 40.140000 12.430000 40.210000 ;
        RECT 12.200000 40.070000 12.500000 40.140000 ;
        RECT 12.270000 40.000000 12.570000 40.070000 ;
        RECT 12.340000 39.930000 12.640000 40.000000 ;
        RECT 12.410000 39.860000 12.710000 39.930000 ;
        RECT 12.480000 39.790000 12.780000 39.860000 ;
        RECT 12.550000 39.720000 12.850000 39.790000 ;
        RECT 12.620000 39.650000 12.920000 39.720000 ;
        RECT 12.690000 39.580000 12.990000 39.650000 ;
        RECT 12.755000  0.000000 13.015000  5.240000 ;
        RECT 12.755000  5.240000 13.015000  5.295000 ;
        RECT 12.755000  5.295000 13.070000  5.350000 ;
        RECT 12.760000 39.510000 13.060000 39.580000 ;
        RECT 12.825000  5.350000 13.125000  5.420000 ;
        RECT 12.830000 39.440000 13.130000 39.510000 ;
        RECT 12.895000  5.420000 13.195000  5.490000 ;
        RECT 12.900000 39.370000 13.200000 39.440000 ;
        RECT 12.965000  5.490000 13.265000  5.560000 ;
        RECT 12.970000 39.300000 13.270000 39.370000 ;
        RECT 13.035000  5.560000 13.335000  5.630000 ;
        RECT 13.040000 39.230000 13.340000 39.300000 ;
        RECT 13.105000  5.630000 13.405000  5.700000 ;
        RECT 13.110000 39.160000 13.410000 39.230000 ;
        RECT 13.175000  5.700000 13.475000  5.770000 ;
        RECT 13.180000 39.090000 13.480000 39.160000 ;
        RECT 13.245000  5.770000 13.545000  5.840000 ;
        RECT 13.250000 39.020000 13.550000 39.090000 ;
        RECT 13.315000  5.840000 13.615000  5.910000 ;
        RECT 13.320000 38.950000 13.620000 39.020000 ;
        RECT 13.385000  5.910000 13.685000  5.980000 ;
        RECT 13.390000 38.880000 13.690000 38.950000 ;
        RECT 13.455000  5.980000 13.755000  6.050000 ;
        RECT 13.460000 38.810000 13.760000 38.880000 ;
        RECT 13.525000  6.050000 13.825000  6.120000 ;
        RECT 13.530000 38.740000 13.830000 38.810000 ;
        RECT 13.595000  6.120000 13.895000  6.190000 ;
        RECT 13.600000 38.670000 13.900000 38.740000 ;
        RECT 13.665000  6.190000 13.965000  6.260000 ;
        RECT 13.670000 38.600000 13.970000 38.670000 ;
        RECT 13.735000  6.260000 14.035000  6.330000 ;
        RECT 13.740000 38.530000 14.040000 38.600000 ;
        RECT 13.805000  6.330000 14.105000  6.400000 ;
        RECT 13.810000 38.460000 14.110000 38.530000 ;
        RECT 13.860000  6.400000 14.175000  6.455000 ;
        RECT 13.880000 38.390000 14.180000 38.460000 ;
        RECT 13.915000  6.455000 14.230000  6.510000 ;
        RECT 13.950000 38.320000 14.250000 38.390000 ;
        RECT 13.970000  6.510000 14.230000  6.565000 ;
        RECT 13.970000  6.565000 14.230000 18.115000 ;
        RECT 13.970000 18.115000 14.230000 18.170000 ;
        RECT 13.970000 18.170000 14.285000 18.225000 ;
        RECT 14.020000 38.250000 14.320000 38.320000 ;
        RECT 14.040000 18.225000 14.340000 18.295000 ;
        RECT 14.090000 38.180000 14.390000 38.250000 ;
        RECT 14.110000 18.295000 14.410000 18.365000 ;
        RECT 14.160000 38.110000 14.460000 38.180000 ;
        RECT 14.180000 18.365000 14.480000 18.435000 ;
        RECT 14.230000 38.040000 14.530000 38.110000 ;
        RECT 14.250000 18.435000 14.550000 18.505000 ;
        RECT 14.300000 37.970000 14.600000 38.040000 ;
        RECT 14.320000 18.505000 14.620000 18.575000 ;
        RECT 14.370000 37.900000 14.670000 37.970000 ;
        RECT 14.390000 18.575000 14.690000 18.645000 ;
        RECT 14.440000 37.830000 14.740000 37.900000 ;
        RECT 14.460000 18.645000 14.760000 18.715000 ;
        RECT 14.510000 37.760000 14.810000 37.830000 ;
        RECT 14.530000 18.715000 14.830000 18.785000 ;
        RECT 14.580000 37.690000 14.880000 37.760000 ;
        RECT 14.600000 18.785000 14.900000 18.855000 ;
        RECT 14.650000 37.620000 14.950000 37.690000 ;
        RECT 14.670000 18.855000 14.970000 18.925000 ;
        RECT 14.720000 37.550000 15.020000 37.620000 ;
        RECT 14.740000 18.925000 15.040000 18.995000 ;
        RECT 14.790000 37.480000 15.090000 37.550000 ;
        RECT 14.810000 18.995000 15.110000 19.065000 ;
        RECT 14.860000 37.410000 15.160000 37.480000 ;
        RECT 14.880000 19.065000 15.180000 19.135000 ;
        RECT 14.915000 37.355000 15.230000 37.410000 ;
        RECT 14.950000 19.135000 15.250000 19.205000 ;
        RECT 14.970000 31.960000 15.285000 32.015000 ;
        RECT 14.970000 32.015000 15.230000 32.070000 ;
        RECT 14.970000 32.070000 15.230000 37.300000 ;
        RECT 14.970000 37.300000 15.230000 37.355000 ;
        RECT 14.995000 31.935000 15.340000 31.960000 ;
        RECT 15.020000 19.205000 15.320000 19.275000 ;
        RECT 15.065000 31.865000 15.365000 31.935000 ;
        RECT 15.090000 19.275000 15.390000 19.345000 ;
        RECT 15.135000 31.795000 15.435000 31.865000 ;
        RECT 15.160000 19.345000 15.460000 19.415000 ;
        RECT 15.205000 31.725000 15.505000 31.795000 ;
        RECT 15.230000 19.415000 15.530000 19.485000 ;
        RECT 15.275000 19.485000 15.600000 19.530000 ;
        RECT 15.275000 31.655000 15.575000 31.725000 ;
        RECT 15.330000 19.530000 15.645000 19.585000 ;
        RECT 15.330000 31.600000 15.645000 31.655000 ;
        RECT 15.385000 19.585000 15.645000 19.640000 ;
        RECT 15.385000 19.640000 15.645000 31.545000 ;
        RECT 15.385000 31.545000 15.645000 31.600000 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    ANTENNAGATEAREA  3.240000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580000 0.000000 78.910000 176.480000 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    ANTENNAGATEAREA  3.120000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.250000 43.835000 11.565000 43.890000 ;
        RECT 11.250000 43.890000 11.510000 43.945000 ;
        RECT 11.250000 43.945000 11.510000 47.275000 ;
        RECT 11.250000 47.275000 11.510000 47.330000 ;
        RECT 11.250000 47.330000 11.565000 47.385000 ;
        RECT 11.270000 43.815000 11.620000 43.835000 ;
        RECT 11.320000 47.385000 11.620000 47.455000 ;
        RECT 11.340000 43.745000 11.640000 43.815000 ;
        RECT 11.390000 47.455000 11.690000 47.525000 ;
        RECT 11.410000 43.675000 11.710000 43.745000 ;
        RECT 11.460000 47.525000 11.760000 47.595000 ;
        RECT 11.480000 43.605000 11.780000 43.675000 ;
        RECT 11.530000 47.595000 11.830000 47.665000 ;
        RECT 11.550000 43.535000 11.850000 43.605000 ;
        RECT 11.600000 47.665000 11.900000 47.735000 ;
        RECT 11.620000 43.465000 11.920000 43.535000 ;
        RECT 11.670000 47.735000 11.970000 47.805000 ;
        RECT 11.680000 47.805000 12.040000 47.815000 ;
        RECT 11.690000 43.395000 11.990000 43.465000 ;
        RECT 11.750000 47.815000 13.850000 47.885000 ;
        RECT 11.760000 43.325000 12.060000 43.395000 ;
        RECT 11.820000 47.885000 13.920000 47.955000 ;
        RECT 11.830000 43.255000 12.130000 43.325000 ;
        RECT 11.890000 47.955000 13.990000 48.025000 ;
        RECT 11.900000 43.185000 12.200000 43.255000 ;
        RECT 11.940000 48.025000 14.060000 48.075000 ;
        RECT 11.970000 43.115000 12.270000 43.185000 ;
        RECT 12.040000 43.045000 12.340000 43.115000 ;
        RECT 12.110000 42.975000 12.410000 43.045000 ;
        RECT 12.180000 42.905000 12.480000 42.975000 ;
        RECT 12.250000 42.835000 12.550000 42.905000 ;
        RECT 12.320000 42.765000 12.620000 42.835000 ;
        RECT 12.390000 42.695000 12.690000 42.765000 ;
        RECT 12.460000 42.625000 12.760000 42.695000 ;
        RECT 12.530000 42.555000 12.830000 42.625000 ;
        RECT 12.600000 42.485000 12.900000 42.555000 ;
        RECT 12.670000 42.415000 12.970000 42.485000 ;
        RECT 12.740000 42.345000 13.040000 42.415000 ;
        RECT 12.810000 42.275000 13.110000 42.345000 ;
        RECT 12.880000 42.205000 13.180000 42.275000 ;
        RECT 12.950000 42.135000 13.250000 42.205000 ;
        RECT 13.020000 42.065000 13.320000 42.135000 ;
        RECT 13.090000 41.995000 13.390000 42.065000 ;
        RECT 13.160000 41.925000 13.460000 41.995000 ;
        RECT 13.230000 41.855000 13.530000 41.925000 ;
        RECT 13.300000 41.785000 13.600000 41.855000 ;
        RECT 13.370000 41.715000 13.670000 41.785000 ;
        RECT 13.440000 41.645000 13.740000 41.715000 ;
        RECT 13.510000 41.575000 13.810000 41.645000 ;
        RECT 13.565000 41.520000 13.880000 41.575000 ;
        RECT 13.620000 40.430000 13.935000 40.485000 ;
        RECT 13.620000 40.485000 13.880000 40.540000 ;
        RECT 13.620000 40.540000 13.880000 41.465000 ;
        RECT 13.620000 41.465000 13.880000 41.520000 ;
        RECT 13.640000 40.410000 13.990000 40.430000 ;
        RECT 13.710000 40.340000 14.010000 40.410000 ;
        RECT 13.780000 40.270000 14.080000 40.340000 ;
        RECT 13.810000 48.075000 14.110000 48.145000 ;
        RECT 13.850000 40.200000 14.150000 40.270000 ;
        RECT 13.880000 48.145000 14.180000 48.215000 ;
        RECT 13.920000 40.130000 14.220000 40.200000 ;
        RECT 13.950000 48.215000 14.250000 48.285000 ;
        RECT 13.990000 40.060000 14.290000 40.130000 ;
        RECT 14.020000 48.285000 14.320000 48.355000 ;
        RECT 14.060000 39.990000 14.360000 40.060000 ;
        RECT 14.090000 48.355000 14.390000 48.425000 ;
        RECT 14.130000 39.920000 14.430000 39.990000 ;
        RECT 14.160000 48.425000 14.460000 48.495000 ;
        RECT 14.180000 39.870000 15.420000 39.920000 ;
        RECT 14.195000 58.050000 14.835000 58.310000 ;
        RECT 14.210000 58.035000 14.820000 58.050000 ;
        RECT 14.230000 48.495000 14.530000 48.565000 ;
        RECT 14.240000 48.565000 14.600000 48.575000 ;
        RECT 14.250000 39.800000 15.470000 39.870000 ;
        RECT 14.280000 57.965000 14.750000 58.035000 ;
        RECT 14.295000 48.575000 14.610000 48.630000 ;
        RECT 14.320000 39.730000 15.540000 39.800000 ;
        RECT 14.350000 48.630000 14.610000 48.685000 ;
        RECT 14.350000 48.685000 14.610000 57.825000 ;
        RECT 14.350000 57.825000 14.610000 57.860000 ;
        RECT 14.350000 57.860000 14.645000 57.895000 ;
        RECT 14.350000 57.895000 14.680000 57.965000 ;
        RECT 14.390000 39.660000 15.610000 39.730000 ;
        RECT 15.365000 39.605000 15.680000 39.660000 ;
        RECT 15.435000 39.535000 15.735000 39.605000 ;
        RECT 15.505000 39.465000 15.805000 39.535000 ;
        RECT 15.575000 39.395000 15.875000 39.465000 ;
        RECT 15.645000 39.325000 15.945000 39.395000 ;
        RECT 15.715000 39.255000 16.015000 39.325000 ;
        RECT 15.785000 39.185000 16.085000 39.255000 ;
        RECT 15.855000 39.115000 16.155000 39.185000 ;
        RECT 15.925000 39.045000 16.225000 39.115000 ;
        RECT 15.995000 38.975000 16.295000 39.045000 ;
        RECT 16.065000 38.905000 16.365000 38.975000 ;
        RECT 16.135000 38.835000 16.435000 38.905000 ;
        RECT 16.205000 38.765000 16.505000 38.835000 ;
        RECT 16.275000 38.695000 16.575000 38.765000 ;
        RECT 16.310000  0.000000 16.570000  2.210000 ;
        RECT 16.310000  2.210000 16.570000  2.265000 ;
        RECT 16.310000  2.265000 16.625000  2.320000 ;
        RECT 16.345000 38.625000 16.645000 38.695000 ;
        RECT 16.365000 31.560000 16.680000 31.615000 ;
        RECT 16.365000 31.615000 16.625000 31.670000 ;
        RECT 16.365000 31.670000 16.625000 34.210000 ;
        RECT 16.365000 34.210000 16.625000 34.265000 ;
        RECT 16.365000 34.265000 16.680000 34.320000 ;
        RECT 16.370000 31.555000 16.735000 31.560000 ;
        RECT 16.380000  2.320000 16.680000  2.390000 ;
        RECT 16.415000 38.555000 16.715000 38.625000 ;
        RECT 16.435000 31.490000 16.740000 31.555000 ;
        RECT 16.435000 34.320000 16.735000 34.390000 ;
        RECT 16.450000  2.390000 16.750000  2.460000 ;
        RECT 16.485000 38.485000 16.785000 38.555000 ;
        RECT 16.500000 31.425000 16.805000 31.490000 ;
        RECT 16.505000 34.390000 16.805000 34.460000 ;
        RECT 16.520000  2.460000 16.820000  2.530000 ;
        RECT 16.555000 31.370000 16.870000 31.425000 ;
        RECT 16.555000 38.415000 16.855000 38.485000 ;
        RECT 16.575000 34.460000 16.875000 34.530000 ;
        RECT 16.590000  2.530000 16.890000  2.600000 ;
        RECT 16.610000  7.160000 16.925000  7.215000 ;
        RECT 16.610000  7.215000 16.870000  7.270000 ;
        RECT 16.610000  7.270000 16.870000 11.540000 ;
        RECT 16.610000 12.475000 16.870000 31.315000 ;
        RECT 16.610000 31.315000 16.870000 31.370000 ;
        RECT 16.615000 12.470000 16.870000 12.475000 ;
        RECT 16.625000 38.345000 16.925000 38.415000 ;
        RECT 16.635000  7.135000 16.980000  7.160000 ;
        RECT 16.645000 34.530000 16.945000 34.600000 ;
        RECT 16.655000 11.540000 16.870000 11.585000 ;
        RECT 16.660000  2.600000 16.960000  2.670000 ;
        RECT 16.660000 12.425000 16.870000 12.470000 ;
        RECT 16.695000 38.275000 16.995000 38.345000 ;
        RECT 16.700000 11.585000 16.870000 11.630000 ;
        RECT 16.705000  7.065000 17.005000  7.135000 ;
        RECT 16.705000 11.630000 16.870000 11.635000 ;
        RECT 16.705000 11.635000 16.870000 12.380000 ;
        RECT 16.705000 12.380000 16.870000 12.425000 ;
        RECT 16.715000 34.600000 17.015000 34.670000 ;
        RECT 16.730000  2.670000 17.030000  2.740000 ;
        RECT 16.765000 38.205000 17.065000 38.275000 ;
        RECT 16.775000  6.995000 17.075000  7.065000 ;
        RECT 16.785000 34.670000 17.085000 34.740000 ;
        RECT 16.800000  2.740000 17.100000  2.810000 ;
        RECT 16.835000 38.135000 17.135000 38.205000 ;
        RECT 16.845000  6.925000 17.145000  6.995000 ;
        RECT 16.855000 34.740000 17.155000 34.810000 ;
        RECT 16.870000  2.810000 17.170000  2.880000 ;
        RECT 16.905000 38.065000 17.205000 38.135000 ;
        RECT 16.915000  6.855000 17.215000  6.925000 ;
        RECT 16.925000 34.810000 17.225000 34.880000 ;
        RECT 16.940000  2.880000 17.240000  2.950000 ;
        RECT 16.975000 37.995000 17.275000 38.065000 ;
        RECT 16.985000  2.950000 17.310000  2.995000 ;
        RECT 16.985000  6.785000 17.285000  6.855000 ;
        RECT 16.995000 34.880000 17.295000 34.950000 ;
        RECT 17.040000  2.995000 17.355000  3.050000 ;
        RECT 17.040000  6.730000 17.355000  6.785000 ;
        RECT 17.045000 37.925000 17.345000 37.995000 ;
        RECT 17.065000 34.950000 17.365000 35.020000 ;
        RECT 17.095000  3.050000 17.355000  3.105000 ;
        RECT 17.095000  3.105000 17.355000  6.675000 ;
        RECT 17.095000  6.675000 17.355000  6.730000 ;
        RECT 17.115000 37.855000 17.415000 37.925000 ;
        RECT 17.135000 35.020000 17.435000 35.090000 ;
        RECT 17.185000 37.785000 17.485000 37.855000 ;
        RECT 17.205000 35.090000 17.505000 35.160000 ;
        RECT 17.255000 37.715000 17.555000 37.785000 ;
        RECT 17.275000 35.160000 17.575000 35.230000 ;
        RECT 17.325000 37.645000 17.625000 37.715000 ;
        RECT 17.345000 35.230000 17.645000 35.300000 ;
        RECT 17.395000 37.575000 17.695000 37.645000 ;
        RECT 17.415000 35.300000 17.715000 35.370000 ;
        RECT 17.465000 35.370000 17.785000 35.420000 ;
        RECT 17.465000 37.505000 17.765000 37.575000 ;
        RECT 17.520000 35.420000 17.835000 35.475000 ;
        RECT 17.520000 37.450000 17.835000 37.505000 ;
        RECT 17.575000 35.475000 17.835000 35.530000 ;
        RECT 17.575000 35.530000 17.835000 37.395000 ;
        RECT 17.575000 37.395000 17.835000 37.450000 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    ANTENNAGATEAREA  1.620000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815000 0.000000 32.075000 3.965000 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600000 0.000000 26.860000 1.695000 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420000 0.000000 5.650000 4.375000 ;
        RECT 5.420000 4.375000 5.650000 4.425000 ;
        RECT 5.420000 4.425000 5.700000 4.475000 ;
        RECT 5.490000 4.475000 5.750000 4.545000 ;
        RECT 5.560000 4.545000 5.820000 4.615000 ;
        RECT 5.630000 4.615000 5.890000 4.685000 ;
        RECT 5.700000 4.685000 5.960000 4.755000 ;
        RECT 5.770000 4.755000 6.030000 4.825000 ;
        RECT 5.840000 4.825000 6.100000 4.895000 ;
        RECT 5.910000 4.895000 6.170000 4.965000 ;
        RECT 5.910000 6.425000 6.550000 6.685000 ;
        RECT 5.980000 4.965000 6.240000 5.035000 ;
        RECT 6.050000 5.035000 6.310000 5.105000 ;
        RECT 6.120000 5.105000 6.380000 5.175000 ;
        RECT 6.180000 6.390000 6.550000 6.425000 ;
        RECT 6.190000 5.175000 6.450000 5.245000 ;
        RECT 6.220000 5.245000 6.520000 5.275000 ;
        RECT 6.250000 6.320000 6.550000 6.390000 ;
        RECT 6.270000 5.275000 6.550000 5.325000 ;
        RECT 6.320000 5.325000 6.550000 5.375000 ;
        RECT 6.320000 5.375000 6.550000 6.250000 ;
        RECT 6.320000 6.250000 6.550000 6.320000 ;
    END
  END IB_MODE_SEL
  PIN IN
    ANTENNAPARTIALMETALSIDEAREA  303.1200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240000 0.000000 79.570000 176.480000 ;
    END
  END IN
  PIN INP_DIS
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245000 0.000000 45.505000 4.980000 ;
        RECT 45.245000 4.980000 45.505000 5.035000 ;
        RECT 45.245000 5.035000 45.560000 5.090000 ;
        RECT 45.315000 5.090000 45.615000 5.160000 ;
        RECT 45.385000 5.160000 45.685000 5.230000 ;
        RECT 45.455000 5.230000 45.755000 5.300000 ;
        RECT 45.525000 5.300000 45.825000 5.370000 ;
        RECT 45.595000 5.370000 45.895000 5.440000 ;
        RECT 45.665000 5.440000 45.965000 5.510000 ;
        RECT 45.735000 5.510000 46.035000 5.580000 ;
        RECT 45.745000 5.580000 46.105000 5.590000 ;
        RECT 45.800000 5.590000 46.115000 5.645000 ;
        RECT 45.855000 5.645000 46.115000 5.700000 ;
        RECT 45.855000 5.700000 46.115000 6.780000 ;
    END
  END INP_DIS
  PIN IN_H
    ANTENNAPARTIALMETALSIDEAREA  291.9480 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400000   0.000000 1.020000 178.235000 ;
        RECT 0.400000 178.235000 1.020000 178.360000 ;
        RECT 0.400000 178.360000 1.145000 178.485000 ;
        RECT 0.550000 178.485000 1.270000 178.635000 ;
        RECT 0.700000 178.635000 1.420000 178.785000 ;
        RECT 0.850000 178.785000 1.570000 178.935000 ;
        RECT 1.000000 178.935000 1.720000 179.085000 ;
        RECT 1.150000 179.085000 1.870000 179.235000 ;
        RECT 1.300000 179.235000 2.020000 179.385000 ;
        RECT 1.450000 179.385000 2.170000 179.535000 ;
        RECT 1.600000 179.535000 2.320000 179.685000 ;
        RECT 1.750000 179.685000 2.470000 179.835000 ;
        RECT 1.900000 179.835000 2.620000 179.985000 ;
        RECT 2.050000 179.985000 2.770000 180.135000 ;
        RECT 2.200000 180.135000 2.920000 180.285000 ;
        RECT 2.350000 180.285000 3.070000 180.435000 ;
        RECT 2.355000 180.435000 3.220000 180.440000 ;
        RECT 2.505000 180.440000 4.565000 180.590000 ;
        RECT 2.655000 180.590000 4.565000 180.740000 ;
        RECT 2.805000 180.740000 4.565000 180.890000 ;
        RECT 2.955000 180.890000 4.565000 181.040000 ;
        RECT 3.085000 181.040000 4.565000 181.170000 ;
    END
  END IN_H
  PIN OE_N
    ANTENNAGATEAREA  1.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375000  0.000000 3.605000  4.375000 ;
        RECT 3.375000  4.375000 3.605000  4.425000 ;
        RECT 3.375000  4.425000 3.655000  4.475000 ;
        RECT 3.445000  4.475000 3.705000  4.545000 ;
        RECT 3.515000  4.545000 3.775000  4.615000 ;
        RECT 3.585000  4.615000 3.845000  4.685000 ;
        RECT 3.655000  4.685000 3.915000  4.755000 ;
        RECT 3.725000  4.755000 3.985000  4.825000 ;
        RECT 3.770000  4.825000 4.055000  4.870000 ;
        RECT 3.840000  4.870000 5.225000  4.940000 ;
        RECT 3.910000  4.940000 5.295000  5.010000 ;
        RECT 3.980000  5.010000 5.365000  5.080000 ;
        RECT 4.000000  5.080000 5.435000  5.100000 ;
        RECT 5.195000  5.100000 5.455000  5.170000 ;
        RECT 5.265000  5.170000 5.525000  5.240000 ;
        RECT 5.300000  5.240000 5.595000  5.275000 ;
        RECT 5.350000  5.275000 5.630000  5.325000 ;
        RECT 5.400000  5.325000 5.630000  5.375000 ;
        RECT 5.400000  5.375000 5.630000  8.250000 ;
        RECT 5.400000  8.250000 5.630000  8.300000 ;
        RECT 5.400000  8.300000 5.680000  8.350000 ;
        RECT 5.470000  8.350000 5.730000  8.420000 ;
        RECT 5.540000  8.420000 5.800000  8.490000 ;
        RECT 5.610000  8.490000 5.870000  8.560000 ;
        RECT 5.680000  8.560000 5.940000  8.630000 ;
        RECT 5.750000  8.630000 6.010000  8.700000 ;
        RECT 5.820000  8.700000 6.080000  8.770000 ;
        RECT 5.890000  8.770000 6.150000  8.840000 ;
        RECT 5.960000  8.840000 6.220000  8.910000 ;
        RECT 5.965000 42.985000 6.225000 43.625000 ;
        RECT 5.970000 42.980000 6.220000 42.985000 ;
        RECT 5.975000 39.420000 6.255000 39.470000 ;
        RECT 5.975000 39.470000 6.205000 39.520000 ;
        RECT 5.975000 39.520000 6.205000 42.965000 ;
        RECT 5.975000 42.965000 6.205000 42.970000 ;
        RECT 5.975000 42.970000 6.210000 42.975000 ;
        RECT 5.975000 42.975000 6.215000 42.980000 ;
        RECT 5.985000 39.410000 6.305000 39.420000 ;
        RECT 6.030000  8.910000 6.290000  8.980000 ;
        RECT 6.055000 39.340000 6.315000 39.410000 ;
        RECT 6.100000  8.980000 6.360000  9.050000 ;
        RECT 6.125000 39.270000 6.385000 39.340000 ;
        RECT 6.170000  9.050000 6.430000  9.120000 ;
        RECT 6.195000 39.200000 6.455000 39.270000 ;
        RECT 6.240000  9.120000 6.500000  9.190000 ;
        RECT 6.265000 39.130000 6.525000 39.200000 ;
        RECT 6.310000  9.190000 6.570000  9.260000 ;
        RECT 6.335000 39.060000 6.595000 39.130000 ;
        RECT 6.380000  9.260000 6.640000  9.330000 ;
        RECT 6.405000 38.990000 6.665000 39.060000 ;
        RECT 6.450000  9.330000 6.710000  9.400000 ;
        RECT 6.475000  9.400000 6.780000  9.425000 ;
        RECT 6.475000 38.920000 6.735000 38.990000 ;
        RECT 6.525000  9.425000 6.805000  9.475000 ;
        RECT 6.525000 38.870000 6.805000 38.920000 ;
        RECT 6.575000  9.475000 6.805000  9.525000 ;
        RECT 6.575000  9.525000 6.805000 38.820000 ;
        RECT 6.575000 38.820000 6.805000 38.870000 ;
    END
  END OE_N
  PIN OUT
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355000  0.000000 22.615000  6.315000 ;
        RECT 22.355000  6.315000 22.615000  6.370000 ;
        RECT 22.355000  6.370000 22.670000  6.425000 ;
        RECT 22.425000  6.425000 22.725000  6.495000 ;
        RECT 22.495000  6.495000 22.795000  6.565000 ;
        RECT 22.565000  6.565000 22.865000  6.635000 ;
        RECT 22.635000  6.635000 22.935000  6.705000 ;
        RECT 22.655000  6.705000 23.005000  6.725000 ;
        RECT 22.710000  6.725000 23.025000  6.780000 ;
        RECT 22.765000  6.780000 23.025000  6.835000 ;
        RECT 22.765000  6.835000 23.025000 14.375000 ;
        RECT 22.765000 14.375000 23.025000 14.430000 ;
        RECT 22.765000 14.430000 23.080000 14.485000 ;
        RECT 22.835000 14.485000 23.135000 14.555000 ;
        RECT 22.905000 14.555000 23.205000 14.625000 ;
        RECT 22.975000 14.625000 23.275000 14.695000 ;
        RECT 23.045000 14.695000 23.345000 14.765000 ;
        RECT 23.095000 38.695000 23.735000 38.955000 ;
        RECT 23.115000 14.765000 23.415000 14.835000 ;
        RECT 23.185000 14.835000 23.485000 14.905000 ;
        RECT 23.255000 14.905000 23.555000 14.975000 ;
        RECT 23.265000 38.625000 23.735000 38.695000 ;
        RECT 23.325000 14.975000 23.625000 15.045000 ;
        RECT 23.335000 38.555000 23.735000 38.625000 ;
        RECT 23.395000 15.045000 23.695000 15.115000 ;
        RECT 23.405000 38.485000 23.735000 38.555000 ;
        RECT 23.465000 15.115000 23.765000 15.185000 ;
        RECT 23.475000 25.180000 23.790000 25.235000 ;
        RECT 23.475000 25.235000 23.735000 25.290000 ;
        RECT 23.475000 25.290000 23.735000 38.415000 ;
        RECT 23.475000 38.415000 23.735000 38.485000 ;
        RECT 23.510000 25.145000 23.845000 25.180000 ;
        RECT 23.535000 15.185000 23.835000 15.255000 ;
        RECT 23.545000 15.255000 23.905000 15.265000 ;
        RECT 23.545000 25.110000 23.880000 25.145000 ;
        RECT 23.600000 15.265000 23.915000 15.320000 ;
        RECT 23.600000 25.055000 23.915000 25.110000 ;
        RECT 23.655000 15.320000 23.915000 15.375000 ;
        RECT 23.655000 15.375000 23.915000 25.000000 ;
        RECT 23.655000 25.000000 23.915000 25.055000 ;
    END
  END OUT
  PIN PAD
    ANTENNAPARTIALMETALSIDEAREA  216.1550 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 32.115000 125.470000 53.655000 147.015000 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    ANTENNAPARTIALMETALSIDEAREA  3.812250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280000 0.000000 76.920000 1.625000 ;
        RECT 76.280000 1.625000 76.920000 1.695000 ;
        RECT 76.280000 1.695000 76.990000 1.765000 ;
        RECT 76.280000 1.765000 77.060000 1.835000 ;
        RECT 76.280000 1.835000 77.130000 1.905000 ;
        RECT 76.280000 1.905000 77.200000 1.975000 ;
        RECT 76.280000 1.975000 77.270000 2.045000 ;
        RECT 76.280000 2.045000 77.340000 2.055000 ;
        RECT 76.350000 2.055000 77.350000 2.125000 ;
        RECT 76.420000 2.125000 77.420000 2.195000 ;
        RECT 76.490000 2.195000 77.490000 2.265000 ;
        RECT 76.560000 2.265000 77.560000 2.335000 ;
        RECT 76.630000 2.335000 77.630000 2.405000 ;
        RECT 76.700000 2.405000 77.700000 2.475000 ;
        RECT 76.770000 2.475000 77.770000 2.545000 ;
        RECT 76.820000 2.545000 77.840000 2.595000 ;
        RECT 76.890000 2.595000 77.890000 2.665000 ;
        RECT 76.960000 2.665000 77.890000 2.735000 ;
        RECT 77.030000 2.735000 77.890000 2.805000 ;
        RECT 77.100000 2.805000 77.890000 2.875000 ;
        RECT 77.150000 2.875000 77.890000 2.925000 ;
        RECT 77.150000 2.925000 77.890000 5.235000 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    ANTENNAPARTIALMETALSIDEAREA  2.618000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275000 0.000000 68.925000 3.960000 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    ANTENNAPARTIALCUTAREA  4.960000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.600000  7.425000 60.560000   7.575000 ;
        RECT 59.600000  7.575000 60.410000   7.725000 ;
        RECT 59.600000  7.725000 60.385000   7.750000 ;
        RECT 59.600000  7.750000 60.385000  10.610000 ;
        RECT 59.600000 10.610000 60.385000  10.760000 ;
        RECT 59.600000 10.760000 60.535000  10.910000 ;
        RECT 59.600000 10.910000 60.685000  10.935000 ;
        RECT 59.655000  7.370000 60.710000   7.425000 ;
        RECT 59.750000 10.935000 60.710000  11.085000 ;
        RECT 59.805000  7.220000 60.765000   7.370000 ;
        RECT 59.900000 11.085000 60.860000  11.235000 ;
        RECT 59.955000  7.070000 60.915000   7.220000 ;
        RECT 59.985000  7.040000 63.890000   7.070000 ;
        RECT 60.050000 11.235000 61.010000  11.385000 ;
        RECT 60.135000  6.890000 63.890000   7.040000 ;
        RECT 60.200000 11.385000 61.160000  11.535000 ;
        RECT 60.285000  6.740000 63.890000   6.890000 ;
        RECT 60.350000 11.535000 61.310000  11.685000 ;
        RECT 60.435000  6.590000 63.890000   6.740000 ;
        RECT 60.500000 11.685000 61.460000  11.835000 ;
        RECT 60.585000  6.440000 63.890000   6.590000 ;
        RECT 60.610000 19.065000 61.570000  19.215000 ;
        RECT 60.610000 19.215000 61.420000  19.365000 ;
        RECT 60.610000 19.365000 61.395000  19.390000 ;
        RECT 60.610000 19.390000 61.395000  47.360000 ;
        RECT 60.650000 11.835000 61.610000  11.985000 ;
        RECT 60.690000 18.985000 61.720000  19.065000 ;
        RECT 60.735000  6.290000 63.890000   6.440000 ;
        RECT 60.800000 11.985000 61.760000  12.135000 ;
        RECT 60.840000 18.835000 61.800000  18.985000 ;
        RECT 60.950000 12.135000 61.910000  12.285000 ;
        RECT 60.990000 18.685000 61.950000  18.835000 ;
        RECT 61.100000 12.285000 62.060000  12.435000 ;
        RECT 61.140000 12.435000 62.210000  12.475000 ;
        RECT 61.140000 18.535000 62.100000  18.685000 ;
        RECT 61.170000 18.505000 62.250000  18.535000 ;
        RECT 61.290000 12.475000 62.250000  12.625000 ;
        RECT 61.320000 18.355000 62.250000  18.505000 ;
        RECT 61.440000 12.625000 62.250000  12.775000 ;
        RECT 61.470000 12.775000 62.250000  12.805000 ;
        RECT 61.470000 12.805000 62.250000  18.205000 ;
        RECT 61.470000 18.205000 62.250000  18.355000 ;
        RECT 61.710000 35.760000 63.070000  35.910000 ;
        RECT 61.710000 35.910000 62.920000  36.060000 ;
        RECT 61.710000 36.060000 62.780000  36.200000 ;
        RECT 61.710000 36.200000 62.780000  73.005000 ;
        RECT 61.710000 73.005000 62.780000  73.155000 ;
        RECT 61.710000 73.155000 62.930000  73.305000 ;
        RECT 61.710000 73.305000 63.080000  73.455000 ;
        RECT 61.710000 73.455000 63.230000  73.605000 ;
        RECT 61.710000 73.605000 63.380000  73.755000 ;
        RECT 61.710000 73.755000 63.530000  73.905000 ;
        RECT 61.710000 73.905000 63.680000  74.055000 ;
        RECT 61.710000 74.055000 63.830000  74.185000 ;
        RECT 61.735000 35.735000 63.220000  35.760000 ;
        RECT 61.750000 74.185000 63.960000  74.225000 ;
        RECT 61.790000 74.225000 64.000000  74.265000 ;
        RECT 61.885000 35.585000 63.245000  35.735000 ;
        RECT 61.940000 74.265000 68.555000  74.415000 ;
        RECT 62.035000 35.435000 63.395000  35.585000 ;
        RECT 62.090000 74.415000 68.705000  74.565000 ;
        RECT 62.185000 35.285000 63.545000  35.435000 ;
        RECT 62.220000  6.155000 63.890000   6.290000 ;
        RECT 62.235000  7.070000 63.890000   7.220000 ;
        RECT 62.240000 74.565000 68.855000  74.715000 ;
        RECT 62.325000 35.145000 63.695000  35.285000 ;
        RECT 62.370000  6.005000 63.890000   6.155000 ;
        RECT 62.385000  7.220000 63.890000   7.370000 ;
        RECT 62.390000 74.715000 69.005000  74.865000 ;
        RECT 62.475000 34.995000 63.695000  35.145000 ;
        RECT 62.520000  5.855000 63.890000   6.005000 ;
        RECT 62.535000  7.370000 63.890000   7.520000 ;
        RECT 62.540000 74.865000 69.155000  75.015000 ;
        RECT 62.625000 17.825000 63.890000  18.070000 ;
        RECT 62.625000 18.070000 63.795000  18.165000 ;
        RECT 62.625000 18.165000 63.700000  18.260000 ;
        RECT 62.625000 18.260000 63.695000  18.265000 ;
        RECT 62.625000 18.265000 63.695000  34.845000 ;
        RECT 62.625000 34.845000 63.695000  34.995000 ;
        RECT 62.630000 17.820000 63.890000  17.825000 ;
        RECT 62.670000  5.705000 63.890000   5.855000 ;
        RECT 62.685000  7.520000 63.890000   7.670000 ;
        RECT 62.690000 75.015000 69.305000  75.165000 ;
        RECT 62.725000 17.725000 63.890000  17.820000 ;
        RECT 62.820000  0.000000 63.890000   5.555000 ;
        RECT 62.820000  5.555000 63.890000   5.705000 ;
        RECT 62.820000  7.670000 63.890000   7.805000 ;
        RECT 62.820000  7.805000 63.890000  17.630000 ;
        RECT 62.820000 17.630000 63.890000  17.725000 ;
        RECT 62.840000 75.165000 69.455000  75.315000 ;
        RECT 62.860000 75.315000 69.605000  75.335000 ;
        RECT 67.870000 75.335000 69.625000  75.400000 ;
        RECT 67.935000 75.400000 69.690000  75.465000 ;
        RECT 67.940000 75.465000 69.755000  75.470000 ;
        RECT 68.090000 75.470000 69.760000  75.620000 ;
        RECT 68.240000 75.620000 69.760000  75.770000 ;
        RECT 68.390000 75.770000 69.760000  75.920000 ;
        RECT 68.540000 75.920000 69.760000  76.070000 ;
        RECT 68.690000 76.070000 69.760000  76.220000 ;
        RECT 68.690000 76.220000 69.760000 101.910000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.000000 106.585000 12.500000 118.955000 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    ANTENNAPARTIALCUTAREA  0.160000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.390000 1.185000 78.210000 1.465000 ;
        RECT 77.470000 1.125000 78.120000 1.185000 ;
        RECT 77.540000 1.055000 78.050000 1.125000 ;
        RECT 77.610000 0.000000 77.870000 0.875000 ;
        RECT 77.610000 0.875000 77.870000 0.930000 ;
        RECT 77.610000 0.930000 77.925000 0.985000 ;
        RECT 77.610000 0.985000 77.980000 1.055000 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    ANTENNAPARTIALMETALSIDEAREA  85.19250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.230000 50.760000 76.475000 50.805000 ;
        RECT 76.230000 50.805000 76.430000 50.850000 ;
        RECT 76.230000 50.850000 76.430000 52.425000 ;
        RECT 76.230000 52.425000 76.430000 52.470000 ;
        RECT 76.230000 52.470000 76.475000 52.515000 ;
        RECT 76.280000 50.710000 76.520000 50.760000 ;
        RECT 76.300000 52.515000 76.520000 52.585000 ;
        RECT 76.350000 50.640000 76.570000 50.710000 ;
        RECT 76.370000 52.585000 76.590000 52.655000 ;
        RECT 76.420000 50.570000 76.640000 50.640000 ;
        RECT 76.440000 52.655000 76.660000 52.725000 ;
        RECT 76.490000 50.500000 76.710000 50.570000 ;
        RECT 76.510000 52.725000 76.730000 52.795000 ;
        RECT 76.560000 50.430000 76.780000 50.500000 ;
        RECT 76.580000 52.795000 76.800000 52.865000 ;
        RECT 76.630000 50.360000 76.850000 50.430000 ;
        RECT 76.650000 52.865000 76.870000 52.935000 ;
        RECT 76.700000 50.290000 76.920000 50.360000 ;
        RECT 76.720000 52.935000 76.940000 53.005000 ;
        RECT 76.770000 50.220000 76.990000 50.290000 ;
        RECT 76.790000 53.005000 77.010000 53.075000 ;
        RECT 76.825000 53.075000 77.080000 53.110000 ;
        RECT 76.840000 50.150000 77.060000 50.220000 ;
        RECT 76.870000 53.110000 77.115000 53.155000 ;
        RECT 76.900000 96.210000 77.130000 96.225000 ;
        RECT 76.910000 50.080000 77.130000 50.150000 ;
        RECT 76.915000 53.155000 77.115000 53.200000 ;
        RECT 76.915000 53.200000 77.115000 96.195000 ;
        RECT 76.915000 96.195000 77.115000 96.210000 ;
        RECT 76.980000 50.010000 77.200000 50.080000 ;
        RECT 77.050000 49.940000 77.270000 50.010000 ;
        RECT 77.120000 49.870000 77.340000 49.940000 ;
        RECT 77.190000 49.800000 77.410000 49.870000 ;
        RECT 77.260000 49.730000 77.480000 49.800000 ;
        RECT 77.330000 49.660000 77.550000 49.730000 ;
        RECT 77.400000 49.590000 77.620000 49.660000 ;
        RECT 77.470000 49.520000 77.690000 49.590000 ;
        RECT 77.540000 49.450000 77.760000 49.520000 ;
        RECT 77.610000 49.380000 77.830000 49.450000 ;
        RECT 77.680000 49.310000 77.900000 49.380000 ;
        RECT 77.750000 49.240000 77.970000 49.310000 ;
        RECT 77.820000 49.170000 78.040000 49.240000 ;
        RECT 77.890000 49.100000 78.110000 49.170000 ;
        RECT 77.960000 49.030000 78.180000 49.100000 ;
        RECT 78.030000 48.960000 78.250000 49.030000 ;
        RECT 78.100000 48.890000 78.320000 48.960000 ;
        RECT 78.170000 48.820000 78.390000 48.890000 ;
        RECT 78.240000 48.750000 78.460000 48.820000 ;
        RECT 78.310000 48.680000 78.530000 48.750000 ;
        RECT 78.380000 48.610000 78.600000 48.680000 ;
        RECT 78.450000 48.540000 78.670000 48.610000 ;
        RECT 78.520000 48.470000 78.740000 48.540000 ;
        RECT 78.590000 48.400000 78.810000 48.470000 ;
        RECT 78.615000 10.265000 78.910000 10.340000 ;
        RECT 78.615000 10.340000 78.860000 10.390000 ;
        RECT 78.615000 10.390000 78.810000 10.440000 ;
        RECT 78.615000 10.440000 78.805000 10.445000 ;
        RECT 78.615000 10.445000 78.805000 16.245000 ;
        RECT 78.615000 16.245000 78.805000 16.285000 ;
        RECT 78.615000 16.285000 78.845000 16.325000 ;
        RECT 78.620000 10.260000 78.910000 10.265000 ;
        RECT 78.660000 48.330000 78.880000 48.400000 ;
        RECT 78.665000 10.215000 78.910000 10.260000 ;
        RECT 78.685000 16.325000 78.885000 16.395000 ;
        RECT 78.705000  0.000000 78.905000  1.125000 ;
        RECT 78.705000  1.125000 78.905000  1.130000 ;
        RECT 78.705000  1.130000 78.910000  1.215000 ;
        RECT 78.710000  1.215000 78.910000  1.220000 ;
        RECT 78.710000  1.220000 78.910000 10.170000 ;
        RECT 78.710000 10.170000 78.910000 10.215000 ;
        RECT 78.730000 48.260000 78.950000 48.330000 ;
        RECT 78.755000 16.395000 78.955000 16.465000 ;
        RECT 78.800000 48.190000 79.020000 48.260000 ;
        RECT 78.825000 16.465000 79.025000 16.535000 ;
        RECT 78.870000 48.120000 79.090000 48.190000 ;
        RECT 78.895000 16.535000 79.095000 16.605000 ;
        RECT 78.940000 48.050000 79.160000 48.120000 ;
        RECT 78.965000 16.605000 79.165000 16.675000 ;
        RECT 79.010000 47.980000 79.230000 48.050000 ;
        RECT 79.035000 16.675000 79.235000 16.745000 ;
        RECT 79.080000 47.910000 79.300000 47.980000 ;
        RECT 79.105000 16.745000 79.305000 16.815000 ;
        RECT 79.150000 47.840000 79.370000 47.910000 ;
        RECT 79.175000 16.815000 79.375000 16.885000 ;
        RECT 79.220000 47.770000 79.440000 47.840000 ;
        RECT 79.240000 16.885000 79.445000 16.950000 ;
        RECT 79.270000 47.720000 79.510000 47.770000 ;
        RECT 79.280000 16.950000 79.510000 16.990000 ;
        RECT 79.320000 16.990000 79.510000 17.030000 ;
        RECT 79.320000 17.030000 79.510000 47.670000 ;
        RECT 79.320000 47.670000 79.510000 47.720000 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    ANTENNAPARTIALMETALSIDEAREA  165.2660 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715000 0.000000 79.915000 96.000000 ;
    END
  END TIE_LO_ESD
  PIN VTRIP_SEL
    ANTENNAGATEAREA  0.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130000 0.000000 6.390000 1.440000 ;
        RECT 6.130000 1.440000 6.390000 1.495000 ;
        RECT 6.130000 1.495000 6.445000 1.550000 ;
        RECT 6.200000 1.550000 6.500000 1.620000 ;
        RECT 6.270000 1.620000 6.570000 1.690000 ;
        RECT 6.340000 1.690000 6.640000 1.760000 ;
        RECT 6.410000 1.760000 6.710000 1.830000 ;
        RECT 6.480000 1.830000 6.780000 1.900000 ;
        RECT 6.550000 1.900000 6.850000 1.970000 ;
        RECT 6.620000 1.970000 6.920000 2.040000 ;
        RECT 6.690000 2.040000 6.990000 2.110000 ;
        RECT 6.760000 2.110000 7.060000 2.180000 ;
        RECT 6.830000 2.180000 7.130000 2.250000 ;
        RECT 6.900000 2.250000 7.200000 2.320000 ;
        RECT 6.970000 2.320000 7.270000 2.390000 ;
        RECT 7.040000 2.390000 7.340000 2.460000 ;
        RECT 7.110000 2.460000 7.410000 2.530000 ;
        RECT 7.180000 2.530000 7.480000 2.600000 ;
        RECT 7.250000 2.600000 7.550000 2.670000 ;
        RECT 7.320000 2.670000 7.620000 2.740000 ;
        RECT 7.390000 2.740000 7.690000 2.810000 ;
        RECT 7.460000 2.810000 7.760000 2.880000 ;
        RECT 7.530000 2.880000 7.830000 2.950000 ;
        RECT 7.600000 2.950000 7.900000 3.020000 ;
        RECT 7.670000 3.020000 7.970000 3.090000 ;
        RECT 7.740000 3.090000 8.040000 3.160000 ;
        RECT 7.810000 3.160000 8.110000 3.230000 ;
        RECT 7.880000 3.230000 8.180000 3.300000 ;
        RECT 7.950000 3.300000 8.250000 3.370000 ;
        RECT 8.020000 3.370000 8.320000 3.440000 ;
        RECT 8.090000 3.440000 8.390000 3.510000 ;
        RECT 8.160000 3.510000 8.460000 3.580000 ;
        RECT 8.230000 3.580000 8.530000 3.650000 ;
        RECT 8.300000 3.650000 8.600000 3.720000 ;
        RECT 8.335000 3.720000 8.670000 3.755000 ;
        RECT 8.390000 3.755000 8.705000 3.810000 ;
        RECT 8.445000 3.810000 8.705000 3.865000 ;
        RECT 8.445000 3.865000 8.705000 6.780000 ;
    END
  END VTRIP_SEL
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 8.885000 1.270000 13.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 8.885000 80.000000 13.535000 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 2.035000 1.270000 7.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 2.035000 80.000000 7.485000 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 14.935000 0.965000 18.385000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.035000 14.935000 80.000000 18.385000 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 19.785000 1.270000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 70.035000 1.270000 95.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 19.785000 80.000000 24.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 70.035000 80.000000 95.000000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 64.085000 1.270000 68.535000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 64.085000 80.000000 68.535000 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 36.735000 1.270000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 47.735000 1.270000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 51.645000 1.270000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 56.405000 1.270000 56.735000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 36.735000 80.000000 40.185000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 47.735000 80.000000 48.065000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 51.645000 80.000000 52.825000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 56.405000 80.000000 56.735000 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 41.585000 1.270000 46.235000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 41.585000 80.000000 46.235000 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 175.785000 1.270000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000000 25.835000 1.270000 30.485000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 175.785000 80.000000 200.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 25.835000 80.000000 30.485000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000000 58.235000 1.270000 62.685000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 58.235000 80.000000 62.685000 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000000 31.885000 1.270000 35.335000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730000 31.885000 80.000000 35.335000 ;
    END
  END VSWITCH
  OBS
    LAYER li1 ;
      RECT -0.115000  95.895000 45.710000  95.955000 ;
      RECT -0.115000  95.955000  4.915000 130.220000 ;
      RECT -0.115000 131.275000  4.915000 140.050000 ;
      RECT -0.115000 140.050000  1.495000 140.150000 ;
      RECT -0.115000 145.155000  1.495000 145.210000 ;
      RECT -0.115000 145.210000  4.915000 170.090000 ;
      RECT -0.085000  93.065000  9.000000  95.255000 ;
      RECT -0.085000  95.255000 45.710000  95.895000 ;
      RECT -0.085000 130.220000  4.915000 130.225000 ;
      RECT -0.085000 130.995000  4.915000 131.275000 ;
      RECT -0.085000 170.090000  4.915000 178.645000 ;
      RECT  0.950000  18.885000  1.310000  19.055000 ;
      RECT  0.980000  21.465000  1.310000  21.635000 ;
      RECT  1.120000  22.325000  1.310000  22.495000 ;
      RECT  1.150000  19.745000  1.310000  19.915000 ;
      RECT  1.150000  20.605000  1.310000  20.775000 ;
      RECT  1.690000  45.545000  4.585000  45.715000 ;
      RECT  2.260000 145.155000  4.700000 145.210000 ;
      RECT  5.875000   5.940000  6.405000   6.465000 ;
      RECT  6.490000  88.950000  9.000000  93.065000 ;
      RECT  7.805000   5.400000 67.100000   6.230000 ;
      RECT  9.300000  32.000000  9.660000  36.750000 ;
      RECT 10.330000  32.000000 10.690000  36.750000 ;
      RECT 11.410000  32.000000 11.665000  37.260000 ;
      RECT 11.940000  31.110000 12.365000  36.765000 ;
      RECT 12.610000  32.000000 13.140000  37.260000 ;
      RECT 13.390000  32.000000 13.920000  36.750000 ;
      RECT 14.170000  32.000000 14.700000  36.750000 ;
      RECT 14.170000  36.750000 14.305000  37.260000 ;
      RECT 14.320000  26.760000 14.500000  29.470000 ;
      RECT 14.320000  29.470000 14.670000  29.570000 ;
      RECT 14.320000  29.570000 14.490000  30.110000 ;
      RECT 14.955000  32.000000 15.485000  37.260000 ;
      RECT 15.105000  26.760000 15.635000  29.690000 ;
      RECT 15.730000  32.000000 16.260000  36.750000 ;
      RECT 15.730000 179.435000 68.925000 179.450000 ;
      RECT 15.730000 179.450000 77.885000 179.980000 ;
      RECT 15.730000 179.980000 68.925000 180.205000 ;
      RECT 15.885000  26.760000 16.415000  29.470000 ;
      RECT 16.510000  32.000000 16.950000  37.260000 ;
      RECT 16.670000  26.760000 17.200000  29.690000 ;
      RECT 17.210000  32.000000 17.650000  36.750000 ;
      RECT 18.035000  26.760000 18.450000  29.470000 ;
      RECT 18.140000  32.060000 18.630000  36.750000 ;
      RECT 19.040000  26.760000 19.455000  29.470000 ;
      RECT 19.050000  32.000000 19.580000  36.750000 ;
      RECT 19.790000  26.760000 20.320000  29.470000 ;
      RECT 20.640000  32.000000 21.170000  36.750000 ;
      RECT 21.690000  26.760000 22.130000  29.470000 ;
      RECT 22.170000  32.000000 22.700000  36.755000 ;
      RECT 23.725000  32.000000 24.255000  36.755000 ;
      RECT 23.800000  26.760000 24.160000  29.470000 ;
      RECT 24.340000  25.580000 26.330000  25.905000 ;
      RECT 24.340000  25.905000 24.835000  29.690000 ;
      RECT 25.015000  26.760000 25.545000  29.470000 ;
      RECT 25.675000  32.250000 26.090000  37.000000 ;
      RECT 25.930000  59.095000 28.100000  60.125000 ;
      RECT 25.935000  57.585000 29.370000  58.865000 ;
      RECT 26.225000  19.595000 26.670000  24.375000 ;
      RECT 26.385000  32.250000 26.865000  37.330000 ;
      RECT 26.390000  26.760000 26.750000  29.690000 ;
      RECT 26.525000  67.105000 29.670000  67.815000 ;
      RECT 26.975000  19.600000 27.420000  24.365000 ;
      RECT 27.045000  32.250000 27.575000  37.000000 ;
      RECT 27.490000  63.970000 29.315000  64.550000 ;
      RECT 27.510000  26.490000 28.090000  30.360000 ;
      RECT 27.675000  68.735000 29.670000  69.445000 ;
      RECT 27.830000  32.245000 28.360000  37.330000 ;
      RECT 28.340000  59.180000 28.510000  59.710000 ;
      RECT 28.605000  32.250000 29.135000  37.005000 ;
      RECT 28.680000  18.995000 29.210000  23.750000 ;
      RECT 28.860000  95.125000 45.710000  95.255000 ;
      RECT 29.035000  56.755000 29.565000  57.285000 ;
      RECT 29.390000  18.965000 30.080000  23.745000 ;
      RECT 29.390000  32.250000 29.920000  37.330000 ;
      RECT 30.165000  32.250000 30.695000  37.000000 ;
      RECT 30.270000  18.995000 30.800000  23.745000 ;
      RECT 30.950000  32.250000 31.375000  37.330000 ;
      RECT 31.660000  32.250000 32.085000  37.005000 ;
      RECT 31.820000  18.995000 32.350000  23.745000 ;
      RECT 32.410000  32.060000 33.070000  36.750000 ;
      RECT 33.500000  31.990000 33.930000  37.080000 ;
      RECT 34.305000  31.975000 34.865000  36.750000 ;
      RECT 35.060000  31.990000 35.490000  37.080000 ;
      RECT 35.865000  31.975000 36.425000  36.750000 ;
      RECT 35.870000  26.885000 36.305000  28.235000 ;
      RECT 36.620000  31.990000 37.050000  37.080000 ;
      RECT 37.425000  31.975000 37.985000  36.750000 ;
      RECT 38.180000  31.990000 38.610000  37.080000 ;
      RECT 38.985000  31.975000 39.545000  36.750000 ;
      RECT 39.270000  26.885000 39.690000  28.235000 ;
      RECT 39.685000  95.955000 45.710000  96.105000 ;
      RECT 39.715000  31.990000 40.090000  36.750000 ;
      RECT 40.580000  32.155000 40.900000  36.710000 ;
      RECT 43.380000  24.850000 43.870000  27.560000 ;
      RECT 43.855000 180.205000 44.500000 180.370000 ;
      RECT 44.200000  33.270000 44.390000  36.510000 ;
      RECT 45.310000  36.340000 46.360000  36.970000 ;
      RECT 49.340000  32.065000 51.760000  32.445000 ;
      RECT 51.105000  32.445000 51.760000  33.690000 ;
      RECT 52.050000  24.855000 52.580000  27.565000 ;
      RECT 53.470000  24.855000 54.000000  27.565000 ;
      RECT 54.870000  24.855000 55.400000  27.565000 ;
      RECT 56.725000 180.205000 57.305000 180.370000 ;
      RECT 59.360000   2.260000 59.720000   3.430000 ;
      RECT 61.115000   5.230000 67.290000   5.345000 ;
      RECT 61.115000   5.345000 67.100000   5.400000 ;
      RECT 61.370000   5.080000 67.290000   5.230000 ;
      RECT 61.560000   4.765000 67.290000   5.080000 ;
      RECT 64.375000   0.250000 66.075000   1.000000 ;
      RECT 65.660000   6.230000 67.100000   9.570000 ;
      RECT 66.390000   9.570000 67.100000   9.575000 ;
      RECT 66.390000   9.575000 69.665000   9.745000 ;
      RECT 66.390000   9.745000 71.650000  10.185000 ;
      RECT 68.290000   1.940000 69.255000   3.960000 ;
      RECT 69.165000 128.445000 79.585000 130.115000 ;
      RECT 69.625000 179.435000 77.885000 179.450000 ;
      RECT 69.625000 179.980000 77.885000 180.205000 ;
      RECT 69.665000  10.185000 71.650000  11.425000 ;
      RECT 72.315000   1.940000 74.335000   4.420000 ;
      RECT 73.080000   8.080000 74.910000   8.830000 ;
      RECT 74.910000   5.170000 76.930000   5.800000 ;
      RECT 74.910000   5.800000 79.430000   7.820000 ;
      RECT 77.195000   3.705000 79.430000   4.420000 ;
      RECT 77.195000   4.420000 77.775000   5.170000 ;
      RECT 77.410000   3.700000 79.430000   3.705000 ;
      RECT 77.410000   7.820000 79.430000   8.080000 ;
      RECT 79.880000  19.485000 80.120000  25.015000 ;
      RECT 79.880000  30.115000 80.120000  35.725000 ;
    LAYER met1 ;
      RECT -0.115000  95.895000  1.495000 130.220000 ;
      RECT -0.115000 131.275000  1.495000 170.090000 ;
      RECT  0.000000   0.000000  5.565000   1.560000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000  5.565000   3.155000 ;
      RECT  0.000000   0.000000 62.290000   2.055000 ;
      RECT  0.000000   1.560000  5.565000   1.565000 ;
      RECT  0.000000   1.565000  5.565000   2.055000 ;
      RECT  0.000000   1.565000 35.575000   1.635000 ;
      RECT  0.000000   1.635000 35.505000   1.705000 ;
      RECT  0.000000   1.705000 35.435000   1.775000 ;
      RECT  0.000000   1.775000 35.365000   1.845000 ;
      RECT  0.000000   1.845000 35.295000   1.915000 ;
      RECT  0.000000   1.915000 35.225000   1.985000 ;
      RECT  0.000000   1.985000 35.155000   2.055000 ;
      RECT  0.000000   2.055000  5.565000   2.875000 ;
      RECT  0.000000   2.055000 80.000000 106.585000 ;
      RECT  0.000000   2.875000 11.260000   3.155000 ;
      RECT  0.000000   3.155000 67.995000   4.240000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   3.155000 67.995000  10.335000 ;
      RECT  0.000000   4.240000 76.885000   5.515000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   4.240000 76.885000  10.335000 ;
      RECT  0.000000   5.515000 80.000000  10.335000 ;
      RECT  0.000000  10.335000  1.340000  11.155000 ;
      RECT  0.000000  11.155000  0.750000  12.425000 ;
      RECT  0.000000  12.425000 80.000000  13.120000 ;
      RECT  0.000000  14.320000 76.495000  23.850000 ;
      RECT  0.000000  14.320000 80.000000  16.455000 ;
      RECT  0.000000  17.275000 78.550000  23.850000 ;
      RECT  0.000000  17.275000 78.550000  29.840000 ;
      RECT  0.000000  17.275000 79.605000  19.205000 ;
      RECT  0.000000  17.275000 79.605000  20.650000 ;
      RECT  0.000000  17.275000 79.605000  20.650000 ;
      RECT  0.000000  19.205000 79.605000  20.650000 ;
      RECT  0.000000  20.650000 78.550000  29.840000 ;
      RECT  0.000000  20.650000 79.535000  20.720000 ;
      RECT  0.000000  20.650000 79.535000  20.720000 ;
      RECT  0.000000  20.720000 79.465000  20.790000 ;
      RECT  0.000000  20.720000 79.465000  20.790000 ;
      RECT  0.000000  20.790000 79.395000  20.860000 ;
      RECT  0.000000  20.790000 79.395000  20.860000 ;
      RECT  0.000000  20.860000 79.325000  20.930000 ;
      RECT  0.000000  20.860000 79.325000  20.930000 ;
      RECT  0.000000  20.930000 79.255000  21.000000 ;
      RECT  0.000000  20.930000 79.255000  21.000000 ;
      RECT  0.000000  21.000000 79.185000  21.070000 ;
      RECT  0.000000  21.000000 79.185000  21.070000 ;
      RECT  0.000000  21.070000 79.160000  21.095000 ;
      RECT  0.000000  21.070000 79.160000  21.095000 ;
      RECT  0.000000  23.405000 79.160000  23.475000 ;
      RECT  0.000000  23.405000 79.160000  23.475000 ;
      RECT  0.000000  23.475000 79.230000  23.545000 ;
      RECT  0.000000  23.475000 79.230000  23.545000 ;
      RECT  0.000000  23.545000 79.300000  23.615000 ;
      RECT  0.000000  23.545000 79.300000  23.615000 ;
      RECT  0.000000  23.615000 79.370000  23.685000 ;
      RECT  0.000000  23.615000 79.370000  23.685000 ;
      RECT  0.000000  23.685000 79.440000  23.755000 ;
      RECT  0.000000  23.685000 79.440000  23.755000 ;
      RECT  0.000000  23.755000 79.510000  23.825000 ;
      RECT  0.000000  23.755000 79.510000  23.825000 ;
      RECT  0.000000  23.825000 79.580000  23.850000 ;
      RECT  0.000000  23.825000 79.580000  23.850000 ;
      RECT  0.000000  23.850000 79.605000  25.295000 ;
      RECT  0.000000  25.295000 78.845000  36.005000 ;
      RECT  0.000000  25.295000 78.845000  42.035000 ;
      RECT  0.000000  25.295000 80.000000  29.840000 ;
      RECT  0.000000  29.840000 78.845000  42.035000 ;
      RECT  0.000000  29.840000 79.605000  31.400000 ;
      RECT  0.000000  31.400000 79.535000  31.470000 ;
      RECT  0.000000  31.400000 79.535000  31.470000 ;
      RECT  0.000000  31.470000 79.465000  31.540000 ;
      RECT  0.000000  31.470000 79.465000  31.540000 ;
      RECT  0.000000  31.540000 79.395000  31.610000 ;
      RECT  0.000000  31.540000 79.395000  31.610000 ;
      RECT  0.000000  31.610000 79.325000  31.680000 ;
      RECT  0.000000  31.610000 79.325000  31.680000 ;
      RECT  0.000000  31.680000 79.280000  31.725000 ;
      RECT  0.000000  31.680000 79.280000  31.725000 ;
      RECT  0.000000  31.725000 78.845000  34.115000 ;
      RECT  0.000000  34.115000 79.280000  34.185000 ;
      RECT  0.000000  34.115000 79.280000  34.185000 ;
      RECT  0.000000  34.185000 79.350000  34.255000 ;
      RECT  0.000000  34.185000 79.350000  34.255000 ;
      RECT  0.000000  34.255000 79.420000  34.325000 ;
      RECT  0.000000  34.255000 79.420000  34.325000 ;
      RECT  0.000000  34.325000 79.490000  34.395000 ;
      RECT  0.000000  34.325000 79.490000  34.395000 ;
      RECT  0.000000  34.395000 79.560000  34.440000 ;
      RECT  0.000000  34.395000 79.560000  34.440000 ;
      RECT  0.000000  34.440000 79.605000  36.005000 ;
      RECT  0.000000  36.005000 80.000000  42.035000 ;
      RECT  0.000000  42.035000 78.635000  42.340000 ;
      RECT  0.000000  42.340000 78.565000  42.410000 ;
      RECT  0.000000  42.340000 78.565000  42.410000 ;
      RECT  0.000000  42.410000 78.495000  42.480000 ;
      RECT  0.000000  42.410000 78.495000  42.480000 ;
      RECT  0.000000  42.480000 78.425000  42.550000 ;
      RECT  0.000000  42.480000 78.425000  42.550000 ;
      RECT  0.000000  42.550000 78.355000  42.620000 ;
      RECT  0.000000  42.550000 78.355000  42.620000 ;
      RECT  0.000000  42.620000 78.285000  42.690000 ;
      RECT  0.000000  42.620000 78.285000  42.690000 ;
      RECT  0.000000  42.690000 78.215000  42.760000 ;
      RECT  0.000000  42.690000 78.215000  42.760000 ;
      RECT  0.000000  42.760000 78.145000  42.830000 ;
      RECT  0.000000  42.760000 78.145000  42.830000 ;
      RECT  0.000000  42.830000 78.075000  42.900000 ;
      RECT  0.000000  42.830000 78.075000  42.900000 ;
      RECT  0.000000  42.900000 78.005000  42.970000 ;
      RECT  0.000000  42.900000 78.005000  42.970000 ;
      RECT  0.000000  42.970000 78.000000  42.975000 ;
      RECT  0.000000  42.970000 78.000000  42.975000 ;
      RECT  0.000000  42.975000 78.635000  43.235000 ;
      RECT  0.000000  43.235000 80.000000  44.355000 ;
      RECT  0.000000  44.355000  1.020000  45.010000 ;
      RECT  0.000000  45.010000  0.965000  45.240000 ;
      RECT  0.000000  45.240000  0.895000  45.310000 ;
      RECT  0.000000  45.310000  0.825000  45.380000 ;
      RECT  0.000000  45.380000  0.755000  45.450000 ;
      RECT  0.000000  45.450000  0.685000  45.520000 ;
      RECT  0.000000  45.520000  0.615000  45.590000 ;
      RECT  0.000000  45.590000  0.545000  45.660000 ;
      RECT  0.000000  45.660000  0.475000  45.730000 ;
      RECT  0.000000  45.730000  0.405000  45.800000 ;
      RECT  0.000000  45.800000  0.335000  45.870000 ;
      RECT  0.000000  45.870000  0.265000  45.940000 ;
      RECT  0.000000  45.940000  0.195000  46.010000 ;
      RECT  0.000000  46.010000  0.125000  46.080000 ;
      RECT  0.000000  46.080000  0.055000  46.150000 ;
      RECT  0.000000  46.445000  0.965000  46.580000 ;
      RECT  0.000000  46.580000  1.050000  47.350000 ;
      RECT  0.000000  47.350000 80.000000  93.020000 ;
      RECT  0.000000  93.020000  1.070000  94.660000 ;
      RECT  0.000000  94.660000 11.550000  94.830000 ;
      RECT  0.000000  94.830000  1.985000  95.615000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 130.500000  4.530000 130.715000 ;
      RECT  0.000000 130.715000  1.980000 130.995000 ;
      RECT  0.000000 170.370000  1.980000 178.680000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 15.445000 198.405000 ;
      RECT  0.000000 178.680000 80.000000 179.140000 ;
      RECT  0.000000 179.140000 15.445000 180.290000 ;
      RECT  0.000000 180.290000 15.490000 200.000000 ;
      RECT  0.000000 180.290000 80.000000 198.405000 ;
      RECT  0.000000 198.405000 15.490000 200.000000 ;
      RECT  0.210000  13.400000  0.470000  14.040000 ;
      RECT  0.475000  46.125000  5.000000  46.165000 ;
      RECT  0.545000  46.055000  5.000000  46.125000 ;
      RECT  0.615000  45.985000  5.000000  46.055000 ;
      RECT  0.685000  45.915000  5.000000  45.985000 ;
      RECT  0.750000  11.155000 76.825000  12.425000 ;
      RECT  0.750000  13.120000 80.000000  16.125000 ;
      RECT  0.755000  45.845000  5.000000  45.915000 ;
      RECT  0.825000  45.775000  5.000000  45.845000 ;
      RECT  0.895000  45.705000  5.000000  45.775000 ;
      RECT  0.965000  45.635000  5.000000  45.705000 ;
      RECT  1.035000  45.565000  5.000000  45.635000 ;
      RECT  1.105000  45.495000  5.000000  45.565000 ;
      RECT  1.175000  45.425000  5.000000  45.495000 ;
      RECT  1.245000  45.290000  5.000000  45.355000 ;
      RECT  1.245000  45.355000  5.000000  45.425000 ;
      RECT  1.245000  46.165000  5.000000  46.300000 ;
      RECT  1.300000  44.635000  1.730000  45.290000 ;
      RECT  1.330000  46.300000  2.790000  47.070000 ;
      RECT  1.350000  93.300000  8.265000  94.380000 ;
      RECT  1.620000  10.615000  4.025000  10.875000 ;
      RECT  1.775000  95.615000  1.985000 106.585000 ;
      RECT  1.775000 118.955000  1.985000 130.500000 ;
      RECT  1.775000 130.995000  1.980000 140.430000 ;
      RECT  1.775000 140.430000 80.000000 144.875000 ;
      RECT  1.775000 144.875000  1.980000 170.370000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  2.010000  44.355000 80.000000  45.010000 ;
      RECT  2.260000 130.995000  4.700000 139.510000 ;
      RECT  2.260000 139.510000  4.855000 140.150000 ;
      RECT  2.260000 145.155000  4.700000 178.400000 ;
      RECT  2.265000  95.110000  8.970000  95.900000 ;
      RECT  2.265000  95.900000  4.250000 130.220000 ;
      RECT  3.070000  46.580000 80.000000  47.350000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  3.070000  46.580000 80.000000  93.020000 ;
      RECT  4.305000   8.145000 80.000000  11.150000 ;
      RECT  4.305000  11.150000 76.825000  11.155000 ;
      RECT  4.530000  96.180000 80.000000 127.980000 ;
      RECT  4.530000 125.130000 70.100000 128.135000 ;
      RECT  4.530000 128.135000 68.825000 130.425000 ;
      RECT  4.530000 130.425000 70.100000 130.500000 ;
      RECT  4.530000 130.500000 80.000000 130.715000 ;
      RECT  4.980000 130.715000 80.000000 139.230000 ;
      RECT  4.980000 144.875000 80.000000 178.680000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  4.980000 144.875000 80.000000 179.140000 ;
      RECT  5.135000 139.230000 80.000000 140.430000 ;
      RECT  5.135000 139.230000 80.000000 144.875000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  46.580000 ;
      RECT  5.280000  43.235000 80.000000  47.350000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  43.235000 80.000000  93.020000 ;
      RECT  5.280000  45.010000 80.000000  46.580000 ;
      RECT  5.565000   0.000000  6.890000   1.560000 ;
      RECT  5.565000   1.560000 22.990000   1.565000 ;
      RECT  5.845000   2.335000 10.120000   2.595000 ;
      RECT  7.170000   0.270000 10.715000   1.280000 ;
      RECT  8.545000  93.020000 11.550000  94.660000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT  9.250000  47.350000 80.000000 127.980000 ;
      RECT 10.400000   2.055000 35.085000   2.125000 ;
      RECT 10.400000   2.125000 35.015000   2.195000 ;
      RECT 10.400000   2.195000 34.945000   2.265000 ;
      RECT 10.400000   2.265000 34.880000   2.330000 ;
      RECT 10.400000   2.330000 13.640000   2.335000 ;
      RECT 10.400000   2.335000 11.260000   2.875000 ;
      RECT 10.995000   0.000000 18.955000   1.560000 ;
      RECT 11.540000   2.615000 35.170000   2.685000 ;
      RECT 11.540000   2.685000 35.100000   2.755000 ;
      RECT 11.540000   2.755000 35.070000   2.785000 ;
      RECT 11.540000   2.785000 18.385000   2.790000 ;
      RECT 11.540000   2.790000 13.990000   2.795000 ;
      RECT 11.540000   2.795000 13.985000   2.800000 ;
      RECT 11.540000   2.800000 12.220000   2.835000 ;
      RECT 11.540000   2.835000 12.185000   2.870000 ;
      RECT 11.540000   2.870000 12.180000   2.875000 ;
      RECT 12.300000   3.150000 67.995000   3.155000 ;
      RECT 12.300000   3.150000 67.995000   3.155000 ;
      RECT 12.310000   3.140000 67.995000   3.150000 ;
      RECT 12.310000   3.140000 67.995000   3.150000 ;
      RECT 12.320000   3.130000 67.995000   3.140000 ;
      RECT 12.320000   3.130000 67.995000   3.140000 ;
      RECT 12.345000   3.105000 59.170000   3.130000 ;
      RECT 12.345000   3.105000 59.170000   3.130000 ;
      RECT 12.370000   3.080000 59.170000   3.105000 ;
      RECT 12.370000   3.080000 59.170000   3.105000 ;
      RECT 13.760000   2.610000 35.240000   2.615000 ;
      RECT 14.105000   3.075000 59.170000   3.080000 ;
      RECT 14.105000   3.075000 59.170000   3.080000 ;
      RECT 14.110000   3.070000 59.170000   3.075000 ;
      RECT 14.110000   3.070000 59.170000   3.075000 ;
      RECT 15.725000 179.420000 77.705000 180.010000 ;
      RECT 15.770000 198.685000 56.715000 199.975000 ;
      RECT 18.505000   3.065000 19.370000   3.070000 ;
      RECT 19.235000   0.270000 21.375000   1.280000 ;
      RECT 19.490000   2.785000 28.955000   2.790000 ;
      RECT 21.655000   0.000000 22.990000   1.560000 ;
      RECT 23.270000   0.275000 26.265000   1.285000 ;
      RECT 26.545000   0.000000 33.120000   1.560000 ;
      RECT 26.545000   1.560000 34.265000   1.565000 ;
      RECT 29.075000   3.065000 30.425000   3.070000 ;
      RECT 29.075000   3.065000 30.425000   3.070000 ;
      RECT 30.545000   2.785000 35.065000   2.790000 ;
      RECT 33.400000   0.270000 37.775000   1.280000 ;
      RECT 34.545000   1.280000 37.775000   1.285000 ;
      RECT 35.055000   2.550000 35.245000   2.610000 ;
      RECT 35.125000   2.480000 35.305000   2.550000 ;
      RECT 35.195000   2.410000 35.375000   2.480000 ;
      RECT 35.205000   3.045000 59.170000   3.070000 ;
      RECT 35.205000   3.045000 59.170000   3.070000 ;
      RECT 35.265000   2.340000 35.445000   2.410000 ;
      RECT 35.275000   2.975000 59.170000   3.045000 ;
      RECT 35.275000   2.975000 59.170000   3.045000 ;
      RECT 35.335000   2.270000 35.515000   2.340000 ;
      RECT 35.345000   2.905000 59.170000   2.975000 ;
      RECT 35.345000   2.905000 59.170000   2.975000 ;
      RECT 35.405000   2.200000 35.585000   2.270000 ;
      RECT 35.415000   2.835000 59.170000   2.905000 ;
      RECT 35.415000   2.835000 59.170000   2.905000 ;
      RECT 35.475000   2.130000 35.655000   2.200000 ;
      RECT 35.485000   2.765000 59.170000   2.835000 ;
      RECT 35.485000   2.765000 59.170000   2.835000 ;
      RECT 35.515000   2.090000 43.035000   2.130000 ;
      RECT 35.555000   2.695000 59.170000   2.765000 ;
      RECT 35.555000   2.695000 59.170000   2.765000 ;
      RECT 35.560000   2.690000 42.990000   2.695000 ;
      RECT 35.560000   2.690000 42.990000   2.695000 ;
      RECT 35.585000   2.020000 42.965000   2.090000 ;
      RECT 35.630000   2.620000 42.920000   2.690000 ;
      RECT 35.630000   2.620000 42.920000   2.690000 ;
      RECT 35.655000   1.950000 42.895000   2.020000 ;
      RECT 35.700000   2.550000 42.850000   2.620000 ;
      RECT 35.700000   2.550000 42.850000   2.620000 ;
      RECT 35.770000   2.480000 42.780000   2.550000 ;
      RECT 35.770000   2.480000 42.780000   2.550000 ;
      RECT 35.840000   2.410000 42.710000   2.480000 ;
      RECT 35.840000   2.410000 42.710000   2.480000 ;
      RECT 38.055000   0.000000 40.785000   1.145000 ;
      RECT 38.055000   1.145000 39.110000   1.670000 ;
      RECT 39.390000   1.425000 43.110000   1.495000 ;
      RECT 39.390000   1.495000 43.180000   1.565000 ;
      RECT 39.390000   1.565000 43.250000   1.635000 ;
      RECT 39.390000   1.635000 43.320000   1.685000 ;
      RECT 41.065000   0.270000 41.935000   1.285000 ;
      RECT 42.215000   0.000000 55.320000   1.145000 ;
      RECT 42.875000   2.130000 43.075000   2.180000 ;
      RECT 42.925000   2.180000 43.125000   2.230000 ;
      RECT 42.930000   2.230000 43.175000   2.235000 ;
      RECT 43.000000   2.235000 51.520000   2.305000 ;
      RECT 43.070000   2.305000 51.520000   2.375000 ;
      RECT 43.110000   1.685000 43.370000   1.755000 ;
      RECT 43.110000   2.375000 51.520000   2.415000 ;
      RECT 43.180000   1.755000 43.440000   1.825000 ;
      RECT 43.200000   1.825000 43.510000   1.845000 ;
      RECT 43.270000   1.145000 62.150000   1.190000 ;
      RECT 43.270000   1.845000 47.840000   1.915000 ;
      RECT 43.315000   1.190000 62.150000   1.235000 ;
      RECT 43.340000   1.915000 47.770000   1.985000 ;
      RECT 43.385000   1.235000 47.725000   1.305000 ;
      RECT 43.410000   1.985000 47.700000   2.055000 ;
      RECT 43.430000   2.055000 47.680000   2.075000 ;
      RECT 43.455000   1.305000 47.655000   1.375000 ;
      RECT 43.525000   1.375000 47.585000   1.445000 ;
      RECT 43.595000   1.445000 47.515000   1.515000 ;
      RECT 43.645000   1.515000 47.465000   1.565000 ;
      RECT 47.630000   1.795000 47.910000   1.845000 ;
      RECT 47.680000   1.745000 47.960000   1.795000 ;
      RECT 47.700000   1.725000 55.040000   1.745000 ;
      RECT 47.770000   1.655000 55.040000   1.725000 ;
      RECT 47.840000   1.585000 55.040000   1.655000 ;
      RECT 47.910000   1.515000 55.040000   1.585000 ;
      RECT 50.840000   2.195000 51.520000   2.235000 ;
      RECT 50.880000   2.155000 51.520000   2.195000 ;
      RECT 51.800000   2.025000 54.525000   2.095000 ;
      RECT 51.800000   2.025000 54.525000   2.095000 ;
      RECT 51.800000   2.095000 54.595000   2.165000 ;
      RECT 51.800000   2.095000 54.595000   2.165000 ;
      RECT 51.800000   2.165000 54.665000   2.235000 ;
      RECT 51.800000   2.165000 54.665000   2.235000 ;
      RECT 51.800000   2.235000 54.735000   2.305000 ;
      RECT 51.800000   2.235000 54.735000   2.305000 ;
      RECT 51.800000   2.305000 54.805000   2.375000 ;
      RECT 51.800000   2.305000 54.805000   2.375000 ;
      RECT 51.800000   2.375000 54.875000   2.445000 ;
      RECT 51.800000   2.375000 54.875000   2.445000 ;
      RECT 51.800000   2.445000 54.945000   2.515000 ;
      RECT 51.800000   2.445000 54.945000   2.515000 ;
      RECT 51.800000   2.515000 55.015000   2.585000 ;
      RECT 51.800000   2.515000 55.015000   2.585000 ;
      RECT 51.800000   2.585000 55.085000   2.655000 ;
      RECT 51.800000   2.585000 55.085000   2.655000 ;
      RECT 51.800000   2.655000 59.170000   2.695000 ;
      RECT 54.655000   1.745000 55.040000   1.760000 ;
      RECT 54.670000   1.760000 55.040000   1.775000 ;
      RECT 54.675000   1.775000 55.040000   1.780000 ;
      RECT 54.745000   1.780000 54.875000   1.850000 ;
      RECT 54.815000   1.850000 54.875000   1.920000 ;
      RECT 55.155000   2.060000 59.170000   2.655000 ;
      RECT 55.320000   0.000000 59.170000   1.145000 ;
      RECT 55.320000   1.145000 59.170000   1.235000 ;
      RECT 55.320000   1.235000 59.170000   1.920000 ;
      RECT 55.320000   1.920000 59.170000   2.060000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 71.715000 200.000000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 180.290000 80.000000 198.420000 ;
      RECT 56.995000 198.405000 80.000000 198.420000 ;
      RECT 56.995000 198.420000 71.715000 200.000000 ;
      RECT 59.170000   0.000000 62.150000   1.145000 ;
      RECT 59.170000   1.235000 62.150000   1.920000 ;
      RECT 59.450000   2.200000 59.710000   2.850000 ;
      RECT 59.990000   1.920000 62.150000   2.195000 ;
      RECT 59.990000   2.195000 67.995000   3.130000 ;
      RECT 62.830000   0.000000 80.000000   2.055000 ;
      RECT 62.970000   0.000000 64.095000   1.190000 ;
      RECT 62.970000   1.190000 67.995000   1.960000 ;
      RECT 62.970000   1.960000 67.995000   2.195000 ;
      RECT 64.375000   0.260000 67.295000   0.910000 ;
      RECT 67.575000   0.000000 69.205000   1.190000 ;
      RECT 67.995000   1.190000 69.205000   1.960000 ;
      RECT 68.275000   2.240000 68.925000   3.960000 ;
      RECT 69.105000 128.415000 80.145000 130.145000 ;
      RECT 69.205000   0.000000 80.000000   1.190000 ;
      RECT 69.205000   1.190000 80.000000   1.960000 ;
      RECT 69.205000   1.960000 80.000000   3.365000 ;
      RECT 69.205000   3.365000 76.885000   4.240000 ;
      RECT 70.380000 128.260000 80.145000 128.415000 ;
      RECT 70.380000 130.145000 80.145000 130.220000 ;
      RECT 71.995000 198.700000 76.855000 200.000000 ;
      RECT 76.775000  16.735000 77.415000  16.995000 ;
      RECT 77.105000  11.430000 77.365000  12.145000 ;
      RECT 77.135000 198.420000 80.000000 200.000000 ;
      RECT 77.165000   3.645000 77.805000   5.235000 ;
      RECT 77.645000  11.150000 80.000000  12.425000 ;
      RECT 77.695000  16.455000 80.000000  17.275000 ;
      RECT 77.985000 179.140000 80.000000 180.290000 ;
      RECT 78.085000   3.365000 80.000000   5.515000 ;
      RECT 78.705000  42.665000 79.175000  42.695000 ;
      RECT 78.775000  42.595000 79.175000  42.665000 ;
      RECT 78.830000  21.375000 80.115000  23.125000 ;
      RECT 78.845000  42.525000 79.175000  42.595000 ;
      RECT 78.915000  42.315000 79.175000  42.455000 ;
      RECT 78.915000  42.455000 79.175000  42.525000 ;
      RECT 78.915000  42.695000 79.175000  42.955000 ;
      RECT 79.125000  32.005000 80.115000  33.835000 ;
      RECT 79.325000  21.325000 80.115000  21.375000 ;
      RECT 79.345000  23.125000 80.115000  23.195000 ;
      RECT 79.395000  21.255000 80.115000  21.325000 ;
      RECT 79.415000  23.195000 80.115000  23.265000 ;
      RECT 79.455000  42.035000 80.000000  43.235000 ;
      RECT 79.465000  21.185000 80.115000  21.255000 ;
      RECT 79.465000  31.935000 80.115000  32.005000 ;
      RECT 79.465000  33.835000 80.115000  33.905000 ;
      RECT 79.485000  23.265000 80.115000  23.335000 ;
      RECT 79.535000  21.115000 80.115000  21.185000 ;
      RECT 79.535000  31.865000 80.115000  31.935000 ;
      RECT 79.535000  33.905000 80.115000  33.975000 ;
      RECT 79.555000  23.335000 80.115000  23.405000 ;
      RECT 79.605000  17.275000 80.000000  19.205000 ;
      RECT 79.605000  21.045000 80.115000  21.115000 ;
      RECT 79.605000  31.795000 80.115000  31.865000 ;
      RECT 79.605000  33.975000 80.115000  34.045000 ;
      RECT 79.625000  23.405000 80.115000  23.475000 ;
      RECT 79.675000  20.975000 80.115000  21.045000 ;
      RECT 79.675000  31.725000 80.115000  31.795000 ;
      RECT 79.675000  34.045000 80.115000  34.115000 ;
      RECT 79.695000  23.475000 80.115000  23.545000 ;
      RECT 79.745000  20.905000 80.115000  20.975000 ;
      RECT 79.745000  31.655000 80.115000  31.725000 ;
      RECT 79.745000  34.115000 80.115000  34.185000 ;
      RECT 79.765000  23.545000 80.115000  23.615000 ;
      RECT 79.815000  20.835000 80.115000  20.905000 ;
      RECT 79.815000  31.585000 80.115000  31.655000 ;
      RECT 79.815000  34.185000 80.115000  34.255000 ;
      RECT 79.835000  23.615000 80.115000  23.685000 ;
      RECT 79.885000  19.485000 80.115000  20.765000 ;
      RECT 79.885000  20.765000 80.115000  20.835000 ;
      RECT 79.885000  23.685000 80.115000  23.735000 ;
      RECT 79.885000  23.735000 80.115000  25.015000 ;
      RECT 79.885000  30.120000 80.115000  31.515000 ;
      RECT 79.885000  31.515000 80.115000  31.585000 ;
      RECT 79.885000  34.255000 80.115000  34.325000 ;
      RECT 79.885000  34.325000 80.115000  35.725000 ;
    LAYER met2 ;
      RECT  0.000000   0.000000  3.095000   4.590000 ;
      RECT  0.000000   0.000000  3.235000   4.535000 ;
      RECT  0.000000   4.535000  3.940000   5.240000 ;
      RECT  0.000000   4.590000  3.095000   4.660000 ;
      RECT  0.000000   4.590000  3.095000   4.660000 ;
      RECT  0.000000   4.660000  3.165000   4.730000 ;
      RECT  0.000000   4.660000  3.165000   4.730000 ;
      RECT  0.000000   4.730000  3.235000   4.800000 ;
      RECT  0.000000   4.730000  3.235000   4.800000 ;
      RECT  0.000000   4.800000  3.305000   4.870000 ;
      RECT  0.000000   4.800000  3.305000   4.870000 ;
      RECT  0.000000   4.870000  3.375000   4.940000 ;
      RECT  0.000000   4.870000  3.375000   4.940000 ;
      RECT  0.000000   4.940000  3.445000   5.010000 ;
      RECT  0.000000   4.940000  3.445000   5.010000 ;
      RECT  0.000000   5.010000  3.515000   5.080000 ;
      RECT  0.000000   5.010000  3.515000   5.080000 ;
      RECT  0.000000   5.080000  3.585000   5.150000 ;
      RECT  0.000000   5.080000  3.585000   5.150000 ;
      RECT  0.000000   5.150000  3.655000   5.220000 ;
      RECT  0.000000   5.150000  3.655000   5.220000 ;
      RECT  0.000000   5.220000  3.725000   5.290000 ;
      RECT  0.000000   5.220000  3.725000   5.290000 ;
      RECT  0.000000   5.240000  5.260000   5.435000 ;
      RECT  0.000000   5.290000  3.795000   5.360000 ;
      RECT  0.000000   5.290000  3.795000   5.360000 ;
      RECT  0.000000   5.360000  3.865000   5.380000 ;
      RECT  0.000000   5.360000  3.865000   5.380000 ;
      RECT  0.000000   5.380000  5.010000   5.435000 ;
      RECT  0.000000   5.380000  5.010000   5.435000 ;
      RECT  0.000000   5.435000  5.065000   5.490000 ;
      RECT  0.000000   5.435000  5.065000   5.490000 ;
      RECT  0.000000   5.435000  5.260000   8.410000 ;
      RECT  0.000000   5.490000  5.120000   8.495000 ;
      RECT  0.000000   8.410000  6.435000   9.585000 ;
      RECT  0.000000   8.465000  5.120000   8.535000 ;
      RECT  0.000000   8.465000  5.120000   8.535000 ;
      RECT  0.000000   8.535000  5.190000   8.605000 ;
      RECT  0.000000   8.535000  5.190000   8.605000 ;
      RECT  0.000000   8.605000  5.260000   8.675000 ;
      RECT  0.000000   8.605000  5.260000   8.675000 ;
      RECT  0.000000   8.675000  5.330000   8.745000 ;
      RECT  0.000000   8.675000  5.330000   8.745000 ;
      RECT  0.000000   8.745000  5.400000   8.815000 ;
      RECT  0.000000   8.745000  5.400000   8.815000 ;
      RECT  0.000000   8.815000  5.470000   8.885000 ;
      RECT  0.000000   8.815000  5.470000   8.885000 ;
      RECT  0.000000   8.885000  5.540000   8.955000 ;
      RECT  0.000000   8.885000  5.540000   8.955000 ;
      RECT  0.000000   8.955000  5.610000   9.025000 ;
      RECT  0.000000   8.955000  5.610000   9.025000 ;
      RECT  0.000000   9.025000  5.680000   9.095000 ;
      RECT  0.000000   9.025000  5.680000   9.095000 ;
      RECT  0.000000   9.095000  5.750000   9.165000 ;
      RECT  0.000000   9.095000  5.750000   9.165000 ;
      RECT  0.000000   9.165000  5.820000   9.235000 ;
      RECT  0.000000   9.165000  5.820000   9.235000 ;
      RECT  0.000000   9.235000  5.890000   9.305000 ;
      RECT  0.000000   9.235000  5.890000   9.305000 ;
      RECT  0.000000   9.305000  5.960000   9.375000 ;
      RECT  0.000000   9.305000  5.960000   9.375000 ;
      RECT  0.000000   9.375000  6.030000   9.445000 ;
      RECT  0.000000   9.375000  6.030000   9.445000 ;
      RECT  0.000000   9.445000  6.100000   9.515000 ;
      RECT  0.000000   9.445000  6.100000   9.515000 ;
      RECT  0.000000   9.515000  6.170000   9.585000 ;
      RECT  0.000000   9.515000  6.170000   9.585000 ;
      RECT  0.000000   9.585000  6.240000   9.640000 ;
      RECT  0.000000   9.585000  6.240000   9.640000 ;
      RECT  0.000000   9.585000  6.435000  38.760000 ;
      RECT  0.000000   9.640000  6.295000  38.705000 ;
      RECT  0.000000  38.705000  6.225000  38.775000 ;
      RECT  0.000000  38.705000  6.225000  38.775000 ;
      RECT  0.000000  38.760000  5.835000  39.360000 ;
      RECT  0.000000  38.775000  6.155000  38.845000 ;
      RECT  0.000000  38.775000  6.155000  38.845000 ;
      RECT  0.000000  38.845000  6.085000  38.915000 ;
      RECT  0.000000  38.845000  6.085000  38.915000 ;
      RECT  0.000000  38.915000  6.015000  38.985000 ;
      RECT  0.000000  38.915000  6.015000  38.985000 ;
      RECT  0.000000  38.985000  5.945000  39.055000 ;
      RECT  0.000000  38.985000  5.945000  39.055000 ;
      RECT  0.000000  39.055000  5.875000  39.125000 ;
      RECT  0.000000  39.055000  5.875000  39.125000 ;
      RECT  0.000000  39.125000  5.805000  39.195000 ;
      RECT  0.000000  39.125000  5.805000  39.195000 ;
      RECT  0.000000  39.195000  5.735000  39.265000 ;
      RECT  0.000000  39.195000  5.735000  39.265000 ;
      RECT  0.000000  39.265000  5.695000  39.305000 ;
      RECT  0.000000  39.265000  5.695000  39.305000 ;
      RECT  0.000000  39.305000  5.685000  53.625000 ;
      RECT  0.000000  39.305000  5.695000  42.860000 ;
      RECT  0.000000  39.360000  5.835000  42.915000 ;
      RECT  0.000000  42.860000  5.690000  42.865000 ;
      RECT  0.000000  42.860000  5.690000  42.865000 ;
      RECT  0.000000  42.865000  5.685000  42.870000 ;
      RECT  0.000000  42.865000  5.685000  42.870000 ;
      RECT  0.000000  42.870000  5.685000  43.905000 ;
      RECT  0.000000  42.915000  5.825000  42.925000 ;
      RECT  0.000000  42.925000  5.825000  43.765000 ;
      RECT  0.000000  43.765000  8.055000  44.015000 ;
      RECT  0.000000  43.905000  7.915000  53.625000 ;
      RECT  0.000000  43.905000  7.945000  43.930000 ;
      RECT  0.000000  43.905000  7.945000  43.930000 ;
      RECT  0.000000  43.930000  7.920000  43.955000 ;
      RECT  0.000000  43.930000  7.920000  43.955000 ;
      RECT  0.000000  43.955000  7.915000  43.960000 ;
      RECT  0.000000  43.955000  7.915000  43.960000 ;
      RECT  0.000000  43.960000  7.915000  53.625000 ;
      RECT  0.000000  44.015000  8.055000  53.680000 ;
      RECT  0.000000  53.625000  7.845000  53.695000 ;
      RECT  0.000000  53.625000  7.845000  53.695000 ;
      RECT  0.000000  53.680000  7.835000  53.900000 ;
      RECT  0.000000  53.695000  7.775000  53.765000 ;
      RECT  0.000000  53.695000  7.775000  53.765000 ;
      RECT  0.000000  53.765000  7.705000  53.835000 ;
      RECT  0.000000  53.765000  7.705000  53.835000 ;
      RECT  0.000000  53.835000  7.695000  53.845000 ;
      RECT  0.000000  53.835000  7.695000  53.845000 ;
      RECT  0.000000  53.845000  7.695000  55.685000 ;
      RECT  0.000000  53.900000  7.835000  55.740000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.035000  73.840000 ;
      RECT  0.000000  55.685000  7.625000  55.755000 ;
      RECT  0.000000  55.685000  7.625000  55.755000 ;
      RECT  0.000000  55.740000  7.175000  56.400000 ;
      RECT  0.000000  55.755000  7.555000  55.825000 ;
      RECT  0.000000  55.755000  7.555000  55.825000 ;
      RECT  0.000000  55.825000  7.485000  55.895000 ;
      RECT  0.000000  55.825000  7.485000  55.895000 ;
      RECT  0.000000  55.895000  7.415000  55.965000 ;
      RECT  0.000000  55.895000  7.415000  55.965000 ;
      RECT  0.000000  55.965000  7.345000  56.035000 ;
      RECT  0.000000  55.965000  7.345000  56.035000 ;
      RECT  0.000000  56.035000  7.275000  56.105000 ;
      RECT  0.000000  56.035000  7.275000  56.105000 ;
      RECT  0.000000  56.105000  7.205000  56.175000 ;
      RECT  0.000000  56.105000  7.205000  56.175000 ;
      RECT  0.000000  56.175000  7.135000  56.245000 ;
      RECT  0.000000  56.175000  7.135000  56.245000 ;
      RECT  0.000000  56.245000  7.065000  56.315000 ;
      RECT  0.000000  56.245000  7.065000  56.315000 ;
      RECT  0.000000  56.315000  7.035000  56.345000 ;
      RECT  0.000000  56.315000  7.035000  56.345000 ;
      RECT  0.000000  56.400000  7.175000  73.785000 ;
      RECT  0.000000  73.785000  7.665000  74.270000 ;
      RECT  0.000000  73.840000  7.035000  73.910000 ;
      RECT  0.000000  73.840000  7.035000  73.910000 ;
      RECT  0.000000  73.910000  7.105000  73.980000 ;
      RECT  0.000000  73.910000  7.105000  73.980000 ;
      RECT  0.000000  73.980000  7.175000  74.050000 ;
      RECT  0.000000  73.980000  7.175000  74.050000 ;
      RECT  0.000000  74.050000  7.245000  74.120000 ;
      RECT  0.000000  74.050000  7.245000  74.120000 ;
      RECT  0.000000  74.120000  7.315000  74.190000 ;
      RECT  0.000000  74.120000  7.315000  74.190000 ;
      RECT  0.000000  74.190000  7.385000  74.260000 ;
      RECT  0.000000  74.190000  7.385000  74.260000 ;
      RECT  0.000000  74.260000  7.455000  74.330000 ;
      RECT  0.000000  74.260000  7.455000  74.330000 ;
      RECT  0.000000  74.270000  7.665000  74.850000 ;
      RECT  0.000000  74.330000  7.525000  74.905000 ;
      RECT  0.000000  74.850000  8.070000  75.255000 ;
      RECT  0.000000  74.905000  7.525000  74.965000 ;
      RECT  0.000000  74.905000  7.525000  74.965000 ;
      RECT  0.000000  74.905000  7.525000  74.975000 ;
      RECT  0.000000  74.965000  7.585000  75.020000 ;
      RECT  0.000000  74.965000  7.585000  75.020000 ;
      RECT  0.000000  74.975000  7.595000  75.045000 ;
      RECT  0.000000  75.020000  7.640000  75.310000 ;
      RECT  0.000000  75.045000  7.665000  75.115000 ;
      RECT  0.000000  75.115000  7.735000  75.185000 ;
      RECT  0.000000  75.185000  7.805000  75.255000 ;
      RECT  0.000000  75.255000  7.875000  75.310000 ;
      RECT  0.000000  75.255000  8.070000  77.055000 ;
      RECT  0.000000  75.310000  7.930000  77.005000 ;
      RECT  0.000000  77.005000  7.640000  78.315000 ;
      RECT  0.000000  77.055000  7.980000  77.145000 ;
      RECT  0.000000  77.145000  7.780000  77.685000 ;
      RECT  0.000000  77.685000 76.775000  96.135000 ;
      RECT  0.000000  77.825000 76.635000  96.080000 ;
      RECT  0.000000  96.080000 76.565000  96.150000 ;
      RECT  0.000000  96.080000 76.565000  96.150000 ;
      RECT  0.000000  96.135000 76.545000  96.365000 ;
      RECT  0.000000  96.150000 76.495000  96.220000 ;
      RECT  0.000000  96.150000 76.495000  96.220000 ;
      RECT  0.000000  96.220000 76.425000  96.290000 ;
      RECT  0.000000  96.220000 76.425000  96.290000 ;
      RECT  0.000000  96.290000 76.355000  96.360000 ;
      RECT  0.000000  96.290000 76.355000  96.360000 ;
      RECT  0.000000  96.360000 76.285000  96.430000 ;
      RECT  0.000000  96.360000 76.285000  96.430000 ;
      RECT  0.000000  96.365000 80.000000 106.585000 ;
      RECT  0.000000  96.430000 76.215000  96.500000 ;
      RECT  0.000000  96.430000 76.215000  96.500000 ;
      RECT  0.000000  96.500000 76.210000  96.505000 ;
      RECT  0.000000  96.500000 76.210000  96.505000 ;
      RECT  0.000000  96.505000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.000000 118.955000 80.000000 200.000000 ;
      RECT  0.740000 106.585000 80.000000 118.955000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT  3.745000   0.000000  5.280000   4.315000 ;
      RECT  3.745000   4.315000  5.280000   4.535000 ;
      RECT  3.885000   0.000000  5.140000   4.260000 ;
      RECT  3.955000   4.260000  5.140000   4.330000 ;
      RECT  3.960000   4.535000  5.475000   4.730000 ;
      RECT  4.025000   4.330000  5.140000   4.400000 ;
      RECT  4.095000   4.400000  5.140000   4.470000 ;
      RECT  4.165000   4.470000  5.140000   4.540000 ;
      RECT  4.215000   4.540000  5.140000   4.590000 ;
      RECT  5.285000   4.730000  5.965000   5.215000 ;
      RECT  5.770000   5.215000  6.180000   5.435000 ;
      RECT  5.770000   5.435000  6.180000   6.190000 ;
      RECT  5.770000   6.190000  6.085000   6.285000 ;
      RECT  5.770000   6.825000  8.305000   6.920000 ;
      RECT  5.770000   6.920000 13.830000   8.190000 ;
      RECT  5.770000   8.190000 13.830000   9.365000 ;
      RECT  5.790000   0.000000  5.990000   1.610000 ;
      RECT  5.790000   1.610000  8.305000   3.925000 ;
      RECT  5.790000   3.925000  8.305000   4.315000 ;
      RECT  5.790000   4.315000  8.305000   5.215000 ;
      RECT  5.845000   2.335000  6.520000   2.405000 ;
      RECT  5.845000   2.405000  6.590000   2.475000 ;
      RECT  5.845000   2.475000  6.660000   2.545000 ;
      RECT  5.845000   2.545000  6.730000   2.595000 ;
      RECT  5.885000   2.595000  6.780000   2.635000 ;
      RECT  5.910000   6.965000  8.165000   7.060000 ;
      RECT  5.910000   7.060000 13.690000   7.345000 ;
      RECT  5.910000   7.345000 13.690000   8.135000 ;
      RECT  5.925000   2.635000  6.820000   2.675000 ;
      RECT  5.930000   1.815000  6.000000   1.885000 ;
      RECT  5.930000   1.885000  6.070000   1.955000 ;
      RECT  5.930000   1.955000  6.140000   2.025000 ;
      RECT  5.930000   2.025000  6.210000   2.095000 ;
      RECT  5.930000   2.095000  6.280000   2.165000 ;
      RECT  5.930000   2.165000  6.350000   2.235000 ;
      RECT  5.930000   2.235000  6.420000   2.305000 ;
      RECT  5.930000   2.305000  6.490000   2.335000 ;
      RECT  5.930000   2.675000  6.860000   2.680000 ;
      RECT  5.930000   2.680000  6.865000   2.750000 ;
      RECT  5.930000   2.750000  6.935000   2.820000 ;
      RECT  5.930000   2.820000  7.005000   2.890000 ;
      RECT  5.930000   2.890000  7.075000   2.960000 ;
      RECT  5.930000   2.960000  7.145000   3.030000 ;
      RECT  5.930000   3.030000  7.215000   3.100000 ;
      RECT  5.930000   3.100000  7.285000   3.170000 ;
      RECT  5.930000   3.170000  7.355000   3.240000 ;
      RECT  5.930000   3.240000  7.425000   3.310000 ;
      RECT  5.930000   3.310000  7.495000   3.380000 ;
      RECT  5.930000   3.380000  7.565000   3.450000 ;
      RECT  5.930000   3.450000  7.635000   3.520000 ;
      RECT  5.930000   3.520000  7.705000   3.590000 ;
      RECT  5.930000   3.590000  7.775000   3.660000 ;
      RECT  5.930000   3.660000  7.845000   3.730000 ;
      RECT  5.930000   3.730000  7.915000   3.800000 ;
      RECT  5.930000   3.800000  7.985000   3.870000 ;
      RECT  5.930000   3.870000  8.055000   3.940000 ;
      RECT  5.930000   3.940000  8.125000   3.980000 ;
      RECT  5.930000   3.980000  8.165000   4.260000 ;
      RECT  5.980000   8.135000 13.690000   8.205000 ;
      RECT  5.980000   8.135000 13.690000   8.205000 ;
      RECT  6.000000   4.260000  8.165000   4.330000 ;
      RECT  6.050000   8.205000 13.690000   8.275000 ;
      RECT  6.050000   8.205000 13.690000   8.275000 ;
      RECT  6.070000   4.330000  8.165000   4.400000 ;
      RECT  6.120000   8.275000 13.690000   8.345000 ;
      RECT  6.120000   8.275000 13.690000   8.345000 ;
      RECT  6.140000   4.400000  8.165000   4.470000 ;
      RECT  6.190000   8.345000 13.690000   8.415000 ;
      RECT  6.190000   8.345000 13.690000   8.415000 ;
      RECT  6.210000   4.470000  8.165000   4.540000 ;
      RECT  6.260000   8.415000 13.690000   8.485000 ;
      RECT  6.260000   8.415000 13.690000   8.485000 ;
      RECT  6.280000   4.540000  8.165000   4.610000 ;
      RECT  6.330000   8.485000 13.690000   8.555000 ;
      RECT  6.330000   8.485000 13.690000   8.555000 ;
      RECT  6.345000  39.580000  9.165000  42.905000 ;
      RECT  6.345000  42.905000  9.145000  42.925000 ;
      RECT  6.350000   4.610000  8.165000   4.680000 ;
      RECT  6.365000  42.925000  8.305000  43.765000 ;
      RECT  6.400000   8.555000 13.690000   8.625000 ;
      RECT  6.400000   8.555000 13.690000   8.625000 ;
      RECT  6.420000   4.680000  8.165000   4.750000 ;
      RECT  6.470000   8.625000 13.690000   8.695000 ;
      RECT  6.470000   8.625000 13.690000   8.695000 ;
      RECT  6.485000  39.635000 12.170000  39.705000 ;
      RECT  6.485000  39.635000 12.170000  39.705000 ;
      RECT  6.485000  39.705000 12.100000  39.775000 ;
      RECT  6.485000  39.705000 12.100000  39.775000 ;
      RECT  6.485000  39.775000 12.030000  39.845000 ;
      RECT  6.485000  39.775000 12.030000  39.845000 ;
      RECT  6.485000  39.845000 11.960000  39.915000 ;
      RECT  6.485000  39.845000 11.960000  39.915000 ;
      RECT  6.485000  39.915000 11.890000  39.985000 ;
      RECT  6.485000  39.915000 11.890000  39.985000 ;
      RECT  6.485000  39.985000 11.820000  40.055000 ;
      RECT  6.485000  39.985000 11.820000  40.055000 ;
      RECT  6.485000  40.055000 11.750000  40.125000 ;
      RECT  6.485000  40.055000 11.750000  40.125000 ;
      RECT  6.485000  40.125000 11.680000  40.195000 ;
      RECT  6.485000  40.125000 11.680000  40.195000 ;
      RECT  6.485000  40.195000 11.610000  40.265000 ;
      RECT  6.485000  40.195000 11.610000  40.265000 ;
      RECT  6.485000  40.265000 11.540000  40.335000 ;
      RECT  6.485000  40.265000 11.540000  40.335000 ;
      RECT  6.485000  40.335000 11.470000  40.405000 ;
      RECT  6.485000  40.335000 11.470000  40.405000 ;
      RECT  6.485000  40.405000 11.400000  40.475000 ;
      RECT  6.485000  40.405000 11.400000  40.475000 ;
      RECT  6.485000  40.475000 11.330000  40.545000 ;
      RECT  6.485000  40.475000 11.330000  40.545000 ;
      RECT  6.485000  40.545000 11.260000  40.615000 ;
      RECT  6.485000  40.545000 11.260000  40.615000 ;
      RECT  6.485000  40.615000 11.190000  40.685000 ;
      RECT  6.485000  40.615000 11.190000  40.685000 ;
      RECT  6.485000  40.685000 11.120000  40.755000 ;
      RECT  6.485000  40.685000 11.120000  40.755000 ;
      RECT  6.485000  40.755000 11.050000  40.825000 ;
      RECT  6.485000  40.755000 11.050000  40.825000 ;
      RECT  6.485000  40.825000 10.980000  40.895000 ;
      RECT  6.485000  40.825000 10.980000  40.895000 ;
      RECT  6.485000  40.895000 10.910000  40.965000 ;
      RECT  6.485000  40.895000 10.910000  40.965000 ;
      RECT  6.485000  40.965000 10.840000  41.035000 ;
      RECT  6.485000  40.965000 10.840000  41.035000 ;
      RECT  6.485000  41.035000 10.770000  41.105000 ;
      RECT  6.485000  41.035000 10.770000  41.105000 ;
      RECT  6.485000  41.105000 10.700000  41.175000 ;
      RECT  6.485000  41.105000 10.700000  41.175000 ;
      RECT  6.485000  41.175000 10.630000  41.245000 ;
      RECT  6.485000  41.175000 10.630000  41.245000 ;
      RECT  6.485000  41.245000 10.560000  41.315000 ;
      RECT  6.485000  41.245000 10.560000  41.315000 ;
      RECT  6.485000  41.315000 10.490000  41.385000 ;
      RECT  6.485000  41.315000 10.490000  41.385000 ;
      RECT  6.485000  41.385000 10.420000  41.455000 ;
      RECT  6.485000  41.385000 10.420000  41.455000 ;
      RECT  6.485000  41.455000 10.350000  41.525000 ;
      RECT  6.485000  41.455000 10.350000  41.525000 ;
      RECT  6.485000  41.525000 10.280000  41.595000 ;
      RECT  6.485000  41.525000 10.280000  41.595000 ;
      RECT  6.485000  41.595000 10.210000  41.665000 ;
      RECT  6.485000  41.595000 10.210000  41.665000 ;
      RECT  6.485000  41.665000 10.140000  41.735000 ;
      RECT  6.485000  41.665000 10.140000  41.735000 ;
      RECT  6.485000  41.735000 10.070000  41.805000 ;
      RECT  6.485000  41.735000 10.070000  41.805000 ;
      RECT  6.485000  41.805000 10.000000  41.875000 ;
      RECT  6.485000  41.805000 10.000000  41.875000 ;
      RECT  6.485000  41.875000  9.930000  41.945000 ;
      RECT  6.485000  41.875000  9.930000  41.945000 ;
      RECT  6.485000  41.945000  9.860000  42.015000 ;
      RECT  6.485000  41.945000  9.860000  42.015000 ;
      RECT  6.485000  42.015000  9.790000  42.085000 ;
      RECT  6.485000  42.015000  9.790000  42.085000 ;
      RECT  6.485000  42.085000  9.720000  42.155000 ;
      RECT  6.485000  42.085000  9.720000  42.155000 ;
      RECT  6.485000  42.155000  9.650000  42.225000 ;
      RECT  6.485000  42.155000  9.650000  42.225000 ;
      RECT  6.485000  42.225000  9.580000  42.295000 ;
      RECT  6.485000  42.225000  9.580000  42.295000 ;
      RECT  6.485000  42.295000  9.510000  42.365000 ;
      RECT  6.485000  42.295000  9.510000  42.365000 ;
      RECT  6.485000  42.365000  9.440000  42.435000 ;
      RECT  6.485000  42.365000  9.440000  42.435000 ;
      RECT  6.485000  42.435000  9.370000  42.505000 ;
      RECT  6.485000  42.435000  9.370000  42.505000 ;
      RECT  6.485000  42.505000  9.300000  42.575000 ;
      RECT  6.485000  42.505000  9.300000  42.575000 ;
      RECT  6.485000  42.575000  9.230000  42.645000 ;
      RECT  6.485000  42.575000  9.230000  42.645000 ;
      RECT  6.485000  42.645000  9.160000  42.715000 ;
      RECT  6.485000  42.645000  9.160000  42.715000 ;
      RECT  6.485000  42.715000  9.090000  42.785000 ;
      RECT  6.485000  42.715000  9.090000  42.785000 ;
      RECT  6.485000  42.785000  9.025000  42.850000 ;
      RECT  6.485000  42.785000  9.025000  42.850000 ;
      RECT  6.490000   4.750000  8.165000   4.820000 ;
      RECT  6.495000  42.850000  9.015000  42.860000 ;
      RECT  6.495000  42.850000  9.015000  42.860000 ;
      RECT  6.505000  42.860000  9.005000  42.870000 ;
      RECT  6.505000  42.860000  9.005000  42.870000 ;
      RECT  6.505000  42.870000  8.935000  42.940000 ;
      RECT  6.505000  42.870000  8.935000  42.940000 ;
      RECT  6.505000  42.940000  8.865000  43.010000 ;
      RECT  6.505000  42.940000  8.865000  43.010000 ;
      RECT  6.505000  43.010000  8.795000  43.080000 ;
      RECT  6.505000  43.010000  8.795000  43.080000 ;
      RECT  6.505000  43.080000  8.725000  43.150000 ;
      RECT  6.505000  43.080000  8.725000  43.150000 ;
      RECT  6.505000  43.150000  8.655000  43.220000 ;
      RECT  6.505000  43.150000  8.655000  43.220000 ;
      RECT  6.505000  43.220000  8.585000  43.290000 ;
      RECT  6.505000  43.220000  8.585000  43.290000 ;
      RECT  6.505000  43.290000  8.515000  43.360000 ;
      RECT  6.505000  43.290000  8.515000  43.360000 ;
      RECT  6.505000  43.360000  8.445000  43.430000 ;
      RECT  6.505000  43.360000  8.445000  43.430000 ;
      RECT  6.505000  43.430000  8.375000  43.500000 ;
      RECT  6.505000  43.430000  8.375000  43.500000 ;
      RECT  6.505000  43.500000  8.305000  43.570000 ;
      RECT  6.505000  43.500000  8.305000  43.570000 ;
      RECT  6.505000  43.570000  8.235000  43.640000 ;
      RECT  6.505000  43.570000  8.235000  43.640000 ;
      RECT  6.505000  43.640000  8.165000  43.710000 ;
      RECT  6.505000  43.640000  8.165000  43.710000 ;
      RECT  6.505000  43.710000  8.095000  43.780000 ;
      RECT  6.505000  43.710000  8.095000  43.780000 ;
      RECT  6.505000  43.780000  8.025000  43.850000 ;
      RECT  6.505000  43.780000  8.025000  43.850000 ;
      RECT  6.505000  43.850000  7.970000  43.905000 ;
      RECT  6.505000  43.850000  7.970000  43.905000 ;
      RECT  6.525000  39.595000 12.240000  39.635000 ;
      RECT  6.525000  39.595000 12.240000  39.635000 ;
      RECT  6.530000   0.000000 12.615000   1.380000 ;
      RECT  6.530000   1.380000 12.615000   3.695000 ;
      RECT  6.540000   8.695000 13.690000   8.765000 ;
      RECT  6.540000   8.695000 13.690000   8.765000 ;
      RECT  6.560000   4.820000  8.165000   4.890000 ;
      RECT  6.595000  39.525000 12.280000  39.595000 ;
      RECT  6.595000  39.525000 12.280000  39.595000 ;
      RECT  6.610000   8.765000 13.690000   8.835000 ;
      RECT  6.610000   8.765000 13.690000   8.835000 ;
      RECT  6.630000   4.890000  8.165000   4.960000 ;
      RECT  6.665000  39.455000 12.350000  39.525000 ;
      RECT  6.665000  39.455000 12.350000  39.525000 ;
      RECT  6.670000   0.000000 12.475000   1.325000 ;
      RECT  6.680000   8.835000 13.690000   8.905000 ;
      RECT  6.680000   8.835000 13.690000   8.905000 ;
      RECT  6.690000   5.215000  8.305000   6.825000 ;
      RECT  6.700000   4.960000  8.165000   5.030000 ;
      RECT  6.735000  39.385000 12.420000  39.455000 ;
      RECT  6.735000  39.385000 12.420000  39.455000 ;
      RECT  6.740000   1.325000 12.475000   1.395000 ;
      RECT  6.740000   1.325000 12.475000   1.395000 ;
      RECT  6.750000   8.905000 13.690000   8.975000 ;
      RECT  6.750000   8.905000 13.690000   8.975000 ;
      RECT  6.770000   5.030000  8.165000   5.100000 ;
      RECT  6.805000  39.315000 12.490000  39.385000 ;
      RECT  6.805000  39.315000 12.490000  39.385000 ;
      RECT  6.810000   1.395000 12.475000   1.465000 ;
      RECT  6.810000   1.395000 12.475000   1.465000 ;
      RECT  6.820000   8.975000 13.690000   9.045000 ;
      RECT  6.820000   8.975000 13.690000   9.045000 ;
      RECT  6.830000   5.100000  8.165000   5.160000 ;
      RECT  6.830000   5.160000  8.165000   6.965000 ;
      RECT  6.875000  39.245000 12.560000  39.315000 ;
      RECT  6.875000  39.245000 12.560000  39.315000 ;
      RECT  6.880000   1.465000 12.475000   1.535000 ;
      RECT  6.880000   1.465000 12.475000   1.535000 ;
      RECT  6.890000   9.045000 13.690000   9.115000 ;
      RECT  6.890000   9.045000 13.690000   9.115000 ;
      RECT  6.945000   9.365000 13.830000  18.285000 ;
      RECT  6.945000  18.285000 15.245000  19.700000 ;
      RECT  6.945000  19.700000 15.245000  31.485000 ;
      RECT  6.945000  31.485000 14.830000  31.900000 ;
      RECT  6.945000  31.900000 14.830000  37.240000 ;
      RECT  6.945000  37.240000 13.095000  38.980000 ;
      RECT  6.945000  38.980000 12.495000  39.580000 ;
      RECT  6.945000  39.175000 12.630000  39.245000 ;
      RECT  6.945000  39.175000 12.630000  39.245000 ;
      RECT  6.950000   1.535000 12.475000   1.605000 ;
      RECT  6.950000   1.535000 12.475000   1.605000 ;
      RECT  6.960000   9.115000 13.690000   9.185000 ;
      RECT  6.960000   9.115000 13.690000   9.185000 ;
      RECT  7.015000  39.105000 12.700000  39.175000 ;
      RECT  7.015000  39.105000 12.700000  39.175000 ;
      RECT  7.020000   1.605000 12.475000   1.675000 ;
      RECT  7.020000   1.605000 12.475000   1.675000 ;
      RECT  7.030000   9.185000 13.690000   9.255000 ;
      RECT  7.030000   9.185000 13.690000   9.255000 ;
      RECT  7.085000   9.255000 13.690000   9.310000 ;
      RECT  7.085000   9.255000 13.690000   9.310000 ;
      RECT  7.085000   9.310000 13.690000  18.340000 ;
      RECT  7.085000  18.340000 13.690000  18.410000 ;
      RECT  7.085000  18.340000 13.690000  18.410000 ;
      RECT  7.085000  18.410000 13.760000  18.480000 ;
      RECT  7.085000  18.410000 13.760000  18.480000 ;
      RECT  7.085000  18.480000 13.830000  18.550000 ;
      RECT  7.085000  18.480000 13.830000  18.550000 ;
      RECT  7.085000  18.550000 13.900000  18.620000 ;
      RECT  7.085000  18.550000 13.900000  18.620000 ;
      RECT  7.085000  18.620000 13.970000  18.690000 ;
      RECT  7.085000  18.620000 13.970000  18.690000 ;
      RECT  7.085000  18.690000 14.040000  18.760000 ;
      RECT  7.085000  18.690000 14.040000  18.760000 ;
      RECT  7.085000  18.760000 14.110000  18.830000 ;
      RECT  7.085000  18.760000 14.110000  18.830000 ;
      RECT  7.085000  18.830000 14.180000  18.900000 ;
      RECT  7.085000  18.830000 14.180000  18.900000 ;
      RECT  7.085000  18.900000 14.250000  18.970000 ;
      RECT  7.085000  18.900000 14.250000  18.970000 ;
      RECT  7.085000  18.970000 14.320000  19.040000 ;
      RECT  7.085000  18.970000 14.320000  19.040000 ;
      RECT  7.085000  19.040000 14.390000  19.110000 ;
      RECT  7.085000  19.040000 14.390000  19.110000 ;
      RECT  7.085000  19.110000 14.460000  19.180000 ;
      RECT  7.085000  19.110000 14.460000  19.180000 ;
      RECT  7.085000  19.180000 14.530000  19.250000 ;
      RECT  7.085000  19.180000 14.530000  19.250000 ;
      RECT  7.085000  19.250000 14.600000  19.320000 ;
      RECT  7.085000  19.250000 14.600000  19.320000 ;
      RECT  7.085000  19.320000 14.670000  19.390000 ;
      RECT  7.085000  19.320000 14.670000  19.390000 ;
      RECT  7.085000  19.390000 14.740000  19.460000 ;
      RECT  7.085000  19.390000 14.740000  19.460000 ;
      RECT  7.085000  19.460000 14.810000  19.530000 ;
      RECT  7.085000  19.460000 14.810000  19.530000 ;
      RECT  7.085000  19.530000 14.880000  19.600000 ;
      RECT  7.085000  19.530000 14.880000  19.600000 ;
      RECT  7.085000  19.600000 14.950000  19.670000 ;
      RECT  7.085000  19.600000 14.950000  19.670000 ;
      RECT  7.085000  19.670000 15.020000  19.740000 ;
      RECT  7.085000  19.670000 15.020000  19.740000 ;
      RECT  7.085000  19.740000 15.090000  19.755000 ;
      RECT  7.085000  19.740000 15.090000  19.755000 ;
      RECT  7.085000  19.755000 15.105000  31.430000 ;
      RECT  7.085000  31.430000 15.035000  31.500000 ;
      RECT  7.085000  31.430000 15.035000  31.500000 ;
      RECT  7.085000  31.500000 14.965000  31.570000 ;
      RECT  7.085000  31.500000 14.965000  31.570000 ;
      RECT  7.085000  31.570000 14.895000  31.640000 ;
      RECT  7.085000  31.570000 14.895000  31.640000 ;
      RECT  7.085000  31.640000 14.825000  31.710000 ;
      RECT  7.085000  31.640000 14.825000  31.710000 ;
      RECT  7.085000  31.710000 14.755000  31.780000 ;
      RECT  7.085000  31.710000 14.755000  31.780000 ;
      RECT  7.085000  31.780000 14.690000  31.845000 ;
      RECT  7.085000  31.780000 14.690000  31.845000 ;
      RECT  7.085000  31.845000 14.690000  37.185000 ;
      RECT  7.085000  37.185000 14.620000  37.255000 ;
      RECT  7.085000  37.185000 14.620000  37.255000 ;
      RECT  7.085000  37.255000 14.550000  37.325000 ;
      RECT  7.085000  37.255000 14.550000  37.325000 ;
      RECT  7.085000  37.325000 14.480000  37.395000 ;
      RECT  7.085000  37.325000 14.480000  37.395000 ;
      RECT  7.085000  37.395000 14.410000  37.465000 ;
      RECT  7.085000  37.395000 14.410000  37.465000 ;
      RECT  7.085000  37.465000 14.340000  37.535000 ;
      RECT  7.085000  37.465000 14.340000  37.535000 ;
      RECT  7.085000  37.535000 14.270000  37.605000 ;
      RECT  7.085000  37.535000 14.270000  37.605000 ;
      RECT  7.085000  37.605000 14.200000  37.675000 ;
      RECT  7.085000  37.605000 14.200000  37.675000 ;
      RECT  7.085000  37.675000 14.130000  37.745000 ;
      RECT  7.085000  37.675000 14.130000  37.745000 ;
      RECT  7.085000  37.745000 14.060000  37.815000 ;
      RECT  7.085000  37.745000 14.060000  37.815000 ;
      RECT  7.085000  37.815000 13.990000  37.885000 ;
      RECT  7.085000  37.815000 13.990000  37.885000 ;
      RECT  7.085000  37.885000 13.920000  37.955000 ;
      RECT  7.085000  37.885000 13.920000  37.955000 ;
      RECT  7.085000  37.955000 13.850000  38.025000 ;
      RECT  7.085000  37.955000 13.850000  38.025000 ;
      RECT  7.085000  38.025000 13.780000  38.095000 ;
      RECT  7.085000  38.025000 13.780000  38.095000 ;
      RECT  7.085000  38.095000 13.710000  38.165000 ;
      RECT  7.085000  38.095000 13.710000  38.165000 ;
      RECT  7.085000  38.165000 13.640000  38.235000 ;
      RECT  7.085000  38.165000 13.640000  38.235000 ;
      RECT  7.085000  38.235000 13.570000  38.305000 ;
      RECT  7.085000  38.235000 13.570000  38.305000 ;
      RECT  7.085000  38.305000 13.500000  38.375000 ;
      RECT  7.085000  38.305000 13.500000  38.375000 ;
      RECT  7.085000  38.375000 13.430000  38.445000 ;
      RECT  7.085000  38.375000 13.430000  38.445000 ;
      RECT  7.085000  38.445000 13.360000  38.515000 ;
      RECT  7.085000  38.445000 13.360000  38.515000 ;
      RECT  7.085000  38.515000 13.290000  38.585000 ;
      RECT  7.085000  38.515000 13.290000  38.585000 ;
      RECT  7.085000  38.585000 13.220000  38.655000 ;
      RECT  7.085000  38.585000 13.220000  38.655000 ;
      RECT  7.085000  38.655000 13.150000  38.725000 ;
      RECT  7.085000  38.655000 13.150000  38.725000 ;
      RECT  7.085000  38.725000 13.080000  38.795000 ;
      RECT  7.085000  38.725000 13.080000  38.795000 ;
      RECT  7.085000  38.795000 13.010000  38.865000 ;
      RECT  7.085000  38.795000 13.010000  38.865000 ;
      RECT  7.085000  38.865000 12.940000  38.935000 ;
      RECT  7.085000  38.865000 12.940000  38.935000 ;
      RECT  7.085000  38.935000 12.870000  39.005000 ;
      RECT  7.085000  38.935000 12.870000  39.005000 ;
      RECT  7.085000  39.005000 12.840000  39.035000 ;
      RECT  7.085000  39.005000 12.840000  39.035000 ;
      RECT  7.085000  39.035000 12.770000  39.105000 ;
      RECT  7.085000  39.035000 12.770000  39.105000 ;
      RECT  7.090000   1.675000 12.475000   1.745000 ;
      RECT  7.090000   1.675000 12.475000   1.745000 ;
      RECT  7.160000   1.745000 12.475000   1.815000 ;
      RECT  7.160000   1.745000 12.475000   1.815000 ;
      RECT  7.230000   1.815000 12.475000   1.885000 ;
      RECT  7.230000   1.815000 12.475000   1.885000 ;
      RECT  7.300000   1.885000 12.475000   1.955000 ;
      RECT  7.300000   1.885000 12.475000   1.955000 ;
      RECT  7.370000   1.955000 12.475000   2.025000 ;
      RECT  7.370000   1.955000 12.475000   2.025000 ;
      RECT  7.440000   2.025000 12.475000   2.095000 ;
      RECT  7.440000   2.025000 12.475000   2.095000 ;
      RECT  7.510000   2.095000 12.475000   2.165000 ;
      RECT  7.510000   2.095000 12.475000   2.165000 ;
      RECT  7.580000   2.165000 12.475000   2.235000 ;
      RECT  7.580000   2.165000 12.475000   2.235000 ;
      RECT  7.650000   2.235000 12.475000   2.305000 ;
      RECT  7.650000   2.235000 12.475000   2.305000 ;
      RECT  7.715000  56.630000 14.210000  57.835000 ;
      RECT  7.715000  57.835000 14.055000  57.990000 ;
      RECT  7.715000  57.990000 14.055000  58.450000 ;
      RECT  7.715000  58.450000 76.775000  73.555000 ;
      RECT  7.715000  73.555000 76.775000  74.045000 ;
      RECT  7.720000   2.305000 12.475000   2.375000 ;
      RECT  7.720000   2.305000 12.475000   2.375000 ;
      RECT  7.790000   2.375000 12.475000   2.445000 ;
      RECT  7.790000   2.375000 12.475000   2.445000 ;
      RECT  7.855000  56.685000 14.070000  57.780000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 13.915000  73.500000 ;
      RECT  7.855000  57.780000 14.000000  57.850000 ;
      RECT  7.855000  57.780000 14.000000  57.850000 ;
      RECT  7.855000  57.850000 13.930000  57.920000 ;
      RECT  7.855000  57.850000 13.930000  57.920000 ;
      RECT  7.855000  57.920000 13.915000  57.935000 ;
      RECT  7.855000  57.920000 13.915000  57.935000 ;
      RECT  7.855000  57.935000 13.915000  58.590000 ;
      RECT  7.855000  58.590000 76.635000  73.500000 ;
      RECT  7.860000   2.445000 12.475000   2.515000 ;
      RECT  7.860000   2.445000 12.475000   2.515000 ;
      RECT  7.885000  56.655000 14.070000  56.685000 ;
      RECT  7.885000  56.655000 14.070000  56.685000 ;
      RECT  7.925000  73.500000 76.635000  73.570000 ;
      RECT  7.925000  73.500000 76.635000  73.570000 ;
      RECT  7.930000   2.515000 12.475000   2.585000 ;
      RECT  7.930000   2.515000 12.475000   2.585000 ;
      RECT  7.955000  56.585000 14.070000  56.655000 ;
      RECT  7.955000  56.585000 14.070000  56.655000 ;
      RECT  7.995000  73.570000 76.635000  73.640000 ;
      RECT  7.995000  73.570000 76.635000  73.640000 ;
      RECT  8.000000   2.585000 12.475000   2.655000 ;
      RECT  8.000000   2.585000 12.475000   2.655000 ;
      RECT  8.025000  56.515000 14.070000  56.585000 ;
      RECT  8.025000  56.515000 14.070000  56.585000 ;
      RECT  8.065000  73.640000 76.635000  73.710000 ;
      RECT  8.065000  73.640000 76.635000  73.710000 ;
      RECT  8.070000   2.655000 12.475000   2.725000 ;
      RECT  8.070000   2.655000 12.475000   2.725000 ;
      RECT  8.095000  56.445000 14.070000  56.515000 ;
      RECT  8.095000  56.445000 14.070000  56.515000 ;
      RECT  8.135000  73.710000 76.635000  73.780000 ;
      RECT  8.135000  73.710000 76.635000  73.780000 ;
      RECT  8.140000   2.725000 12.475000   2.795000 ;
      RECT  8.140000   2.725000 12.475000   2.795000 ;
      RECT  8.165000  56.375000 14.070000  56.445000 ;
      RECT  8.165000  56.375000 14.070000  56.445000 ;
      RECT  8.205000  73.780000 76.635000  73.850000 ;
      RECT  8.205000  73.780000 76.635000  73.850000 ;
      RECT  8.205000  74.045000 76.775000  74.620000 ;
      RECT  8.205000  74.620000 76.775000  75.025000 ;
      RECT  8.210000   2.795000 12.475000   2.865000 ;
      RECT  8.210000   2.795000 12.475000   2.865000 ;
      RECT  8.235000  56.305000 14.070000  56.375000 ;
      RECT  8.235000  56.305000 14.070000  56.375000 ;
      RECT  8.275000  73.850000 76.635000  73.920000 ;
      RECT  8.275000  73.850000 76.635000  73.920000 ;
      RECT  8.280000   2.865000 12.475000   2.935000 ;
      RECT  8.280000   2.865000 12.475000   2.935000 ;
      RECT  8.305000  56.235000 14.070000  56.305000 ;
      RECT  8.305000  56.235000 14.070000  56.305000 ;
      RECT  8.345000  73.920000 76.635000  73.990000 ;
      RECT  8.345000  73.920000 76.635000  73.990000 ;
      RECT  8.345000  73.990000 76.635000  74.565000 ;
      RECT  8.350000   2.935000 12.475000   3.005000 ;
      RECT  8.350000   2.935000 12.475000   3.005000 ;
      RECT  8.375000  54.130000 14.210000  55.970000 ;
      RECT  8.375000  55.970000 14.210000  56.630000 ;
      RECT  8.375000  56.165000 14.070000  56.235000 ;
      RECT  8.375000  56.165000 14.070000  56.235000 ;
      RECT  8.415000  74.565000 76.635000  74.635000 ;
      RECT  8.415000  74.565000 76.635000  74.635000 ;
      RECT  8.420000   3.005000 12.475000   3.075000 ;
      RECT  8.420000   3.005000 12.475000   3.075000 ;
      RECT  8.445000  56.095000 14.070000  56.165000 ;
      RECT  8.445000  56.095000 14.070000  56.165000 ;
      RECT  8.485000  74.635000 76.635000  74.705000 ;
      RECT  8.485000  74.635000 76.635000  74.705000 ;
      RECT  8.490000   3.075000 12.475000   3.145000 ;
      RECT  8.490000   3.075000 12.475000   3.145000 ;
      RECT  8.515000  54.185000 14.070000  56.025000 ;
      RECT  8.515000  56.025000 14.070000  56.095000 ;
      RECT  8.515000  56.025000 14.070000  56.095000 ;
      RECT  8.525000  54.175000 14.070000  54.185000 ;
      RECT  8.525000  54.175000 14.070000  54.185000 ;
      RECT  8.555000  74.705000 76.635000  74.775000 ;
      RECT  8.555000  74.705000 76.635000  74.775000 ;
      RECT  8.560000   3.145000 12.475000   3.215000 ;
      RECT  8.560000   3.145000 12.475000   3.215000 ;
      RECT  8.595000  44.245000 11.110000  47.445000 ;
      RECT  8.595000  47.445000 11.880000  48.215000 ;
      RECT  8.595000  48.215000 14.210000  48.745000 ;
      RECT  8.595000  48.745000 14.210000  53.910000 ;
      RECT  8.595000  53.910000 14.210000  54.130000 ;
      RECT  8.595000  54.105000 14.070000  54.175000 ;
      RECT  8.595000  54.105000 14.070000  54.175000 ;
      RECT  8.610000  75.025000 76.775000  77.135000 ;
      RECT  8.610000  77.135000 76.775000  77.225000 ;
      RECT  8.625000  74.775000 76.635000  74.845000 ;
      RECT  8.625000  74.775000 76.635000  74.845000 ;
      RECT  8.630000   3.215000 12.475000   3.285000 ;
      RECT  8.630000   3.215000 12.475000   3.285000 ;
      RECT  8.665000  54.035000 14.070000  54.105000 ;
      RECT  8.665000  54.035000 14.070000  54.105000 ;
      RECT  8.695000  74.845000 76.635000  74.915000 ;
      RECT  8.695000  74.845000 76.635000  74.915000 ;
      RECT  8.700000   3.285000 12.475000   3.355000 ;
      RECT  8.700000   3.285000 12.475000   3.355000 ;
      RECT  8.700000  77.225000 76.775000  77.685000 ;
      RECT  8.735000  44.300000 10.970000  45.265000 ;
      RECT  8.735000  45.335000  8.805000  45.405000 ;
      RECT  8.735000  45.335000  8.805000  45.405000 ;
      RECT  8.735000  45.405000  8.875000  45.475000 ;
      RECT  8.735000  45.405000  8.875000  45.475000 ;
      RECT  8.735000  45.475000  8.945000  45.545000 ;
      RECT  8.735000  45.475000  8.945000  45.545000 ;
      RECT  8.735000  45.545000  9.015000  45.615000 ;
      RECT  8.735000  45.545000  9.015000  45.615000 ;
      RECT  8.735000  45.615000  9.085000  45.685000 ;
      RECT  8.735000  45.615000  9.085000  45.685000 ;
      RECT  8.735000  45.685000  9.155000  45.755000 ;
      RECT  8.735000  45.685000  9.155000  45.755000 ;
      RECT  8.735000  45.755000  9.225000  45.825000 ;
      RECT  8.735000  45.755000  9.225000  45.825000 ;
      RECT  8.735000  45.825000  9.295000  45.895000 ;
      RECT  8.735000  45.825000  9.295000  45.895000 ;
      RECT  8.735000  45.895000  9.365000  45.965000 ;
      RECT  8.735000  45.895000  9.365000  45.965000 ;
      RECT  8.735000  45.965000  9.435000  46.035000 ;
      RECT  8.735000  45.965000  9.435000  46.035000 ;
      RECT  8.735000  46.035000  9.505000  46.105000 ;
      RECT  8.735000  46.035000  9.505000  46.105000 ;
      RECT  8.735000  46.105000  9.575000  46.175000 ;
      RECT  8.735000  46.105000  9.575000  46.175000 ;
      RECT  8.735000  46.175000  9.645000  46.245000 ;
      RECT  8.735000  46.175000  9.645000  46.245000 ;
      RECT  8.735000  46.245000  9.715000  46.315000 ;
      RECT  8.735000  46.245000  9.715000  46.315000 ;
      RECT  8.735000  46.315000  9.785000  46.385000 ;
      RECT  8.735000  46.315000  9.785000  46.385000 ;
      RECT  8.735000  46.385000  9.855000  46.455000 ;
      RECT  8.735000  46.385000  9.855000  46.455000 ;
      RECT  8.735000  46.455000  9.925000  46.525000 ;
      RECT  8.735000  46.455000  9.925000  46.525000 ;
      RECT  8.735000  46.525000  9.995000  46.595000 ;
      RECT  8.735000  46.525000  9.995000  46.595000 ;
      RECT  8.735000  46.595000 10.065000  46.665000 ;
      RECT  8.735000  46.595000 10.065000  46.665000 ;
      RECT  8.735000  46.665000 10.135000  46.735000 ;
      RECT  8.735000  46.665000 10.135000  46.735000 ;
      RECT  8.735000  46.735000 10.205000  46.805000 ;
      RECT  8.735000  46.735000 10.205000  46.805000 ;
      RECT  8.735000  46.805000 10.275000  46.875000 ;
      RECT  8.735000  46.805000 10.275000  46.875000 ;
      RECT  8.735000  46.875000 10.345000  46.945000 ;
      RECT  8.735000  46.875000 10.345000  46.945000 ;
      RECT  8.735000  46.945000 10.415000  47.015000 ;
      RECT  8.735000  46.945000 10.415000  47.015000 ;
      RECT  8.735000  47.015000 10.485000  47.085000 ;
      RECT  8.735000  47.015000 10.485000  47.085000 ;
      RECT  8.735000  47.085000 10.555000  47.155000 ;
      RECT  8.735000  47.085000 10.555000  47.155000 ;
      RECT  8.735000  47.155000 10.625000  47.225000 ;
      RECT  8.735000  47.155000 10.625000  47.225000 ;
      RECT  8.735000  47.225000 10.695000  47.295000 ;
      RECT  8.735000  47.225000 10.695000  47.295000 ;
      RECT  8.735000  47.295000 10.765000  47.365000 ;
      RECT  8.735000  47.295000 10.765000  47.365000 ;
      RECT  8.735000  47.365000 10.835000  47.435000 ;
      RECT  8.735000  47.365000 10.835000  47.435000 ;
      RECT  8.735000  47.435000 10.905000  47.500000 ;
      RECT  8.735000  47.435000 10.905000  47.500000 ;
      RECT  8.735000  47.500000 10.970000  47.570000 ;
      RECT  8.735000  47.500000 10.970000  47.570000 ;
      RECT  8.735000  47.570000 11.040000  47.640000 ;
      RECT  8.735000  47.570000 11.040000  47.640000 ;
      RECT  8.735000  47.640000 11.110000  47.710000 ;
      RECT  8.735000  47.640000 11.110000  47.710000 ;
      RECT  8.735000  47.710000 11.180000  47.780000 ;
      RECT  8.735000  47.710000 11.180000  47.780000 ;
      RECT  8.735000  47.780000 11.250000  47.850000 ;
      RECT  8.735000  47.780000 11.250000  47.850000 ;
      RECT  8.735000  47.850000 11.320000  47.920000 ;
      RECT  8.735000  47.850000 11.320000  47.920000 ;
      RECT  8.735000  47.920000 11.390000  47.990000 ;
      RECT  8.735000  47.920000 11.390000  47.990000 ;
      RECT  8.735000  47.990000 11.460000  48.060000 ;
      RECT  8.735000  47.990000 11.460000  48.060000 ;
      RECT  8.735000  48.060000 11.530000  48.130000 ;
      RECT  8.735000  48.060000 11.530000  48.130000 ;
      RECT  8.735000  48.130000 11.600000  48.200000 ;
      RECT  8.735000  48.130000 11.600000  48.200000 ;
      RECT  8.735000  48.200000 11.670000  48.270000 ;
      RECT  8.735000  48.200000 11.670000  48.270000 ;
      RECT  8.735000  48.270000 11.740000  48.340000 ;
      RECT  8.735000  48.270000 11.740000  48.340000 ;
      RECT  8.735000  48.340000 11.810000  48.355000 ;
      RECT  8.735000  48.340000 11.810000  48.355000 ;
      RECT  8.735000  48.355000 13.625000  48.425000 ;
      RECT  8.735000  48.355000 13.625000  48.425000 ;
      RECT  8.735000  48.425000 13.695000  48.495000 ;
      RECT  8.735000  48.425000 13.695000  48.495000 ;
      RECT  8.735000  48.495000 13.765000  48.565000 ;
      RECT  8.735000  48.495000 13.765000  48.565000 ;
      RECT  8.735000  48.565000 13.835000  48.635000 ;
      RECT  8.735000  48.565000 13.835000  48.635000 ;
      RECT  8.735000  48.635000 13.905000  48.705000 ;
      RECT  8.735000  48.635000 13.905000  48.705000 ;
      RECT  8.735000  48.705000 13.975000  48.775000 ;
      RECT  8.735000  48.705000 13.975000  48.775000 ;
      RECT  8.735000  48.775000 14.045000  48.800000 ;
      RECT  8.735000  48.775000 14.045000  48.800000 ;
      RECT  8.735000  48.800000 14.070000  53.965000 ;
      RECT  8.735000  48.800000 14.070000  56.025000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  48.800000 14.070000  56.685000 ;
      RECT  8.735000  53.965000 14.070000  54.035000 ;
      RECT  8.735000  53.965000 14.070000  54.035000 ;
      RECT  8.750000  74.915000 76.635000  74.970000 ;
      RECT  8.750000  74.915000 76.635000  74.970000 ;
      RECT  8.750000  74.970000 76.635000  77.080000 ;
      RECT  8.755000  44.280000 10.970000  44.300000 ;
      RECT  8.770000   3.355000 12.475000   3.425000 ;
      RECT  8.770000   3.355000 12.475000   3.425000 ;
      RECT  8.795000  77.080000 76.635000  77.125000 ;
      RECT  8.795000  77.080000 76.635000  77.125000 ;
      RECT  8.825000  44.210000 10.970000  44.280000 ;
      RECT  8.840000   3.425000 12.475000   3.495000 ;
      RECT  8.840000   3.425000 12.475000   3.495000 ;
      RECT  8.840000  74.970000 76.635000  96.080000 ;
      RECT  8.840000  74.970000 76.635000  96.080000 ;
      RECT  8.840000  77.125000 76.635000  77.170000 ;
      RECT  8.840000  77.125000 76.635000  77.170000 ;
      RECT  8.845000   3.695000 12.615000   5.410000 ;
      RECT  8.845000   5.410000 13.830000   6.625000 ;
      RECT  8.845000   6.625000 13.830000   6.920000 ;
      RECT  8.895000  44.140000 10.970000  44.210000 ;
      RECT  8.910000   3.495000 12.475000   3.565000 ;
      RECT  8.910000   3.495000 12.475000   3.565000 ;
      RECT  8.965000  44.070000 10.970000  44.140000 ;
      RECT  8.980000   3.565000 12.475000   3.635000 ;
      RECT  8.980000   3.565000 12.475000   3.635000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   1.325000 12.475000   5.465000 ;
      RECT  8.985000   3.635000 12.475000   3.640000 ;
      RECT  8.985000   3.635000 12.475000   3.640000 ;
      RECT  8.985000   5.465000 12.475000   5.535000 ;
      RECT  8.985000   5.465000 12.475000   5.535000 ;
      RECT  8.985000   5.535000 12.545000   5.605000 ;
      RECT  8.985000   5.535000 12.545000   5.605000 ;
      RECT  8.985000   5.605000 12.615000   5.675000 ;
      RECT  8.985000   5.605000 12.615000   5.675000 ;
      RECT  8.985000   5.675000 12.685000   5.745000 ;
      RECT  8.985000   5.675000 12.685000   5.745000 ;
      RECT  8.985000   5.745000 12.755000   5.815000 ;
      RECT  8.985000   5.745000 12.755000   5.815000 ;
      RECT  8.985000   5.815000 12.825000   5.885000 ;
      RECT  8.985000   5.815000 12.825000   5.885000 ;
      RECT  8.985000   5.885000 12.895000   5.955000 ;
      RECT  8.985000   5.885000 12.895000   5.955000 ;
      RECT  8.985000   5.955000 12.965000   6.025000 ;
      RECT  8.985000   5.955000 12.965000   6.025000 ;
      RECT  8.985000   6.025000 13.035000   6.095000 ;
      RECT  8.985000   6.025000 13.035000   6.095000 ;
      RECT  8.985000   6.095000 13.105000   6.165000 ;
      RECT  8.985000   6.095000 13.105000   6.165000 ;
      RECT  8.985000   6.165000 13.175000   6.235000 ;
      RECT  8.985000   6.165000 13.175000   6.235000 ;
      RECT  8.985000   6.235000 13.245000   6.305000 ;
      RECT  8.985000   6.235000 13.245000   6.305000 ;
      RECT  8.985000   6.305000 13.315000   6.375000 ;
      RECT  8.985000   6.305000 13.315000   6.375000 ;
      RECT  8.985000   6.375000 13.385000   6.445000 ;
      RECT  8.985000   6.375000 13.385000   6.445000 ;
      RECT  8.985000   6.445000 13.455000   6.515000 ;
      RECT  8.985000   6.445000 13.455000   6.515000 ;
      RECT  8.985000   6.515000 13.525000   6.585000 ;
      RECT  8.985000   6.515000 13.525000   6.585000 ;
      RECT  8.985000   6.585000 13.595000   6.655000 ;
      RECT  8.985000   6.585000 13.595000   6.655000 ;
      RECT  8.985000   6.655000 13.665000   6.680000 ;
      RECT  8.985000   6.655000 13.665000   6.680000 ;
      RECT  8.985000   6.680000 13.690000   7.060000 ;
      RECT  9.035000  44.000000 10.970000  44.070000 ;
      RECT  9.060000  43.775000 11.110000  44.245000 ;
      RECT  9.105000  43.930000 10.970000  44.000000 ;
      RECT  9.175000  43.860000 10.970000  43.930000 ;
      RECT  9.245000  43.790000 10.970000  43.860000 ;
      RECT  9.315000  43.720000 10.970000  43.790000 ;
      RECT  9.375000  43.660000 10.970000  43.720000 ;
      RECT  9.445000  43.590000 11.030000  43.660000 ;
      RECT  9.515000  43.520000 11.100000  43.590000 ;
      RECT  9.585000  43.450000 11.170000  43.520000 ;
      RECT  9.655000  43.380000 11.240000  43.450000 ;
      RECT  9.725000  43.310000 11.310000  43.380000 ;
      RECT  9.795000  43.240000 11.380000  43.310000 ;
      RECT  9.865000  43.170000 11.450000  43.240000 ;
      RECT  9.935000  43.100000 11.520000  43.170000 ;
      RECT 10.005000  43.030000 11.590000  43.100000 ;
      RECT 10.075000  42.960000 11.660000  43.030000 ;
      RECT 10.145000  42.890000 11.730000  42.960000 ;
      RECT 10.215000  42.820000 11.800000  42.890000 ;
      RECT 10.285000  42.750000 11.870000  42.820000 ;
      RECT 10.355000  42.680000 11.940000  42.750000 ;
      RECT 10.425000  42.610000 12.010000  42.680000 ;
      RECT 10.495000  42.540000 12.080000  42.610000 ;
      RECT 10.565000  42.470000 12.150000  42.540000 ;
      RECT 10.635000  42.400000 12.220000  42.470000 ;
      RECT 10.705000  42.330000 12.290000  42.400000 ;
      RECT 10.775000  42.260000 12.360000  42.330000 ;
      RECT 10.845000  42.190000 12.430000  42.260000 ;
      RECT 10.915000  42.120000 12.500000  42.190000 ;
      RECT 10.985000  42.050000 12.570000  42.120000 ;
      RECT 11.055000  41.980000 12.640000  42.050000 ;
      RECT 11.125000  41.910000 12.710000  41.980000 ;
      RECT 11.195000  41.840000 12.780000  41.910000 ;
      RECT 11.265000  41.770000 12.850000  41.840000 ;
      RECT 11.335000  41.700000 12.920000  41.770000 ;
      RECT 11.405000  41.630000 12.990000  41.700000 ;
      RECT 11.475000  41.560000 13.060000  41.630000 ;
      RECT 11.545000  41.490000 13.130000  41.560000 ;
      RECT 11.615000  41.420000 13.200000  41.490000 ;
      RECT 11.650000  44.005000 29.985000  47.215000 ;
      RECT 11.650000  47.215000 29.985000  47.675000 ;
      RECT 11.685000  41.350000 13.270000  41.420000 ;
      RECT 11.740000  41.295000 13.340000  41.350000 ;
      RECT 11.790000  44.060000 29.845000  47.160000 ;
      RECT 11.810000  41.225000 13.340000  41.295000 ;
      RECT 11.850000  44.000000 29.845000  44.060000 ;
      RECT 11.850000  44.000000 29.845000  44.060000 ;
      RECT 11.860000  47.160000 29.845000  47.230000 ;
      RECT 11.860000  47.160000 29.845000  47.230000 ;
      RECT 11.880000  41.155000 13.340000  41.225000 ;
      RECT 11.920000  43.930000 29.845000  44.000000 ;
      RECT 11.920000  43.930000 29.845000  44.000000 ;
      RECT 11.930000  47.230000 29.845000  47.300000 ;
      RECT 11.930000  47.230000 29.845000  47.300000 ;
      RECT 11.950000  41.085000 13.340000  41.155000 ;
      RECT 11.990000  43.860000 29.845000  43.930000 ;
      RECT 11.990000  43.860000 29.845000  43.930000 ;
      RECT 12.000000  47.300000 29.845000  47.370000 ;
      RECT 12.000000  47.300000 29.845000  47.370000 ;
      RECT 12.020000  41.015000 13.340000  41.085000 ;
      RECT 12.060000  43.790000 29.845000  43.860000 ;
      RECT 12.060000  43.790000 29.845000  43.860000 ;
      RECT 12.070000  47.370000 29.845000  47.440000 ;
      RECT 12.070000  47.370000 29.845000  47.440000 ;
      RECT 12.090000  40.945000 13.340000  41.015000 ;
      RECT 12.130000  43.720000 29.845000  43.790000 ;
      RECT 12.130000  43.720000 29.845000  43.790000 ;
      RECT 12.140000  47.440000 29.845000  47.510000 ;
      RECT 12.140000  47.440000 29.845000  47.510000 ;
      RECT 12.160000  40.875000 13.340000  40.945000 ;
      RECT 12.165000  47.510000 29.845000  47.535000 ;
      RECT 12.165000  47.510000 29.845000  47.535000 ;
      RECT 12.200000  43.650000 29.845000  43.720000 ;
      RECT 12.200000  43.650000 29.845000  43.720000 ;
      RECT 12.230000  40.805000 13.340000  40.875000 ;
      RECT 12.270000  43.580000 29.845000  43.650000 ;
      RECT 12.270000  43.580000 29.845000  43.650000 ;
      RECT 12.300000  40.735000 13.340000  40.805000 ;
      RECT 12.340000  43.510000 29.845000  43.580000 ;
      RECT 12.340000  43.510000 29.845000  43.580000 ;
      RECT 12.370000  40.665000 13.340000  40.735000 ;
      RECT 12.410000  43.440000 29.845000  43.510000 ;
      RECT 12.410000  43.440000 29.845000  43.510000 ;
      RECT 12.440000  40.595000 13.340000  40.665000 ;
      RECT 12.465000  40.370000 13.480000  41.405000 ;
      RECT 12.480000  43.370000 29.845000  43.440000 ;
      RECT 12.480000  43.370000 29.845000  43.440000 ;
      RECT 12.510000  40.525000 13.340000  40.595000 ;
      RECT 12.550000  43.300000 29.845000  43.370000 ;
      RECT 12.550000  43.300000 29.845000  43.370000 ;
      RECT 12.580000  40.455000 13.340000  40.525000 ;
      RECT 12.620000  43.230000 29.845000  43.300000 ;
      RECT 12.620000  43.230000 29.845000  43.300000 ;
      RECT 12.650000  40.385000 13.340000  40.455000 ;
      RECT 12.690000  43.160000 29.845000  43.230000 ;
      RECT 12.690000  43.160000 29.845000  43.230000 ;
      RECT 12.720000  40.315000 13.340000  40.385000 ;
      RECT 12.745000  40.290000 13.340000  40.315000 ;
      RECT 12.760000  43.090000 29.845000  43.160000 ;
      RECT 12.760000  43.090000 29.845000  43.160000 ;
      RECT 12.815000  40.220000 13.365000  40.290000 ;
      RECT 12.830000  43.020000 29.845000  43.090000 ;
      RECT 12.830000  43.020000 29.845000  43.090000 ;
      RECT 12.885000  40.150000 13.435000  40.220000 ;
      RECT 12.900000  42.950000 29.845000  43.020000 ;
      RECT 12.900000  42.950000 29.845000  43.020000 ;
      RECT 12.955000  40.080000 13.505000  40.150000 ;
      RECT 12.970000  42.880000 29.845000  42.950000 ;
      RECT 12.970000  42.880000 29.845000  42.950000 ;
      RECT 13.025000  40.010000 13.575000  40.080000 ;
      RECT 13.040000  42.810000 29.845000  42.880000 ;
      RECT 13.040000  42.810000 29.845000  42.880000 ;
      RECT 13.095000  39.940000 13.645000  40.010000 ;
      RECT 13.110000  42.740000 29.845000  42.810000 ;
      RECT 13.110000  42.740000 29.845000  42.810000 ;
      RECT 13.155000   0.000000 16.170000   2.380000 ;
      RECT 13.155000   2.380000 16.955000   3.160000 ;
      RECT 13.155000   3.160000 16.955000   5.180000 ;
      RECT 13.155000   5.180000 16.955000   6.395000 ;
      RECT 13.165000  39.870000 13.715000  39.940000 ;
      RECT 13.180000  42.670000 29.845000  42.740000 ;
      RECT 13.180000  42.670000 29.845000  42.740000 ;
      RECT 13.235000  39.800000 13.785000  39.870000 ;
      RECT 13.250000  42.600000 29.845000  42.670000 ;
      RECT 13.250000  42.600000 29.845000  42.670000 ;
      RECT 13.295000   0.000000 13.595000   0.070000 ;
      RECT 13.295000   0.000000 13.595000   0.070000 ;
      RECT 13.295000   0.070000 13.665000   0.140000 ;
      RECT 13.295000   0.070000 13.665000   0.140000 ;
      RECT 13.295000   0.140000 13.735000   0.210000 ;
      RECT 13.295000   0.140000 13.735000   0.210000 ;
      RECT 13.295000   0.210000 13.805000   0.280000 ;
      RECT 13.295000   0.210000 13.805000   0.280000 ;
      RECT 13.295000   0.280000 13.875000   0.350000 ;
      RECT 13.295000   0.280000 13.875000   0.350000 ;
      RECT 13.295000   0.350000 13.945000   0.420000 ;
      RECT 13.295000   0.350000 13.945000   0.420000 ;
      RECT 13.295000   0.420000 14.015000   0.490000 ;
      RECT 13.295000   0.420000 14.015000   0.490000 ;
      RECT 13.295000   0.490000 14.085000   0.560000 ;
      RECT 13.295000   0.490000 14.085000   0.560000 ;
      RECT 13.295000   0.560000 14.155000   0.630000 ;
      RECT 13.295000   0.560000 14.155000   0.630000 ;
      RECT 13.295000   0.630000 14.225000   0.700000 ;
      RECT 13.295000   0.630000 14.225000   0.700000 ;
      RECT 13.295000   0.700000 14.295000   0.770000 ;
      RECT 13.295000   0.700000 14.295000   0.770000 ;
      RECT 13.295000   0.770000 14.365000   0.840000 ;
      RECT 13.295000   0.770000 14.365000   0.840000 ;
      RECT 13.295000   0.840000 14.435000   0.910000 ;
      RECT 13.295000   0.840000 14.435000   0.910000 ;
      RECT 13.295000   0.910000 14.505000   0.980000 ;
      RECT 13.295000   0.910000 14.505000   0.980000 ;
      RECT 13.295000   0.980000 14.575000   1.050000 ;
      RECT 13.295000   0.980000 14.575000   1.050000 ;
      RECT 13.295000   1.050000 14.645000   1.120000 ;
      RECT 13.295000   1.050000 14.645000   1.120000 ;
      RECT 13.295000   1.120000 14.715000   1.190000 ;
      RECT 13.295000   1.120000 14.715000   1.190000 ;
      RECT 13.295000   1.190000 14.785000   1.260000 ;
      RECT 13.295000   1.190000 14.785000   1.260000 ;
      RECT 13.295000   1.260000 14.855000   1.330000 ;
      RECT 13.295000   1.260000 14.855000   1.330000 ;
      RECT 13.295000   1.330000 14.925000   1.400000 ;
      RECT 13.295000   1.330000 14.925000   1.400000 ;
      RECT 13.295000   1.400000 14.995000   1.470000 ;
      RECT 13.295000   1.400000 14.995000   1.470000 ;
      RECT 13.295000   1.470000 15.065000   1.540000 ;
      RECT 13.295000   1.470000 15.065000   1.540000 ;
      RECT 13.295000   1.540000 15.135000   1.610000 ;
      RECT 13.295000   1.540000 15.135000   1.610000 ;
      RECT 13.295000   1.610000 15.205000   1.680000 ;
      RECT 13.295000   1.610000 15.205000   1.680000 ;
      RECT 13.295000   1.680000 15.275000   1.750000 ;
      RECT 13.295000   1.680000 15.275000   1.750000 ;
      RECT 13.295000   1.750000 15.345000   1.820000 ;
      RECT 13.295000   1.750000 15.345000   1.820000 ;
      RECT 13.295000   1.820000 15.415000   1.890000 ;
      RECT 13.295000   1.820000 15.415000   1.890000 ;
      RECT 13.295000   1.890000 15.485000   1.960000 ;
      RECT 13.295000   1.890000 15.485000   1.960000 ;
      RECT 13.295000   1.960000 15.555000   2.030000 ;
      RECT 13.295000   1.960000 15.555000   2.030000 ;
      RECT 13.295000   2.030000 15.625000   2.100000 ;
      RECT 13.295000   2.030000 15.625000   2.100000 ;
      RECT 13.295000   2.100000 15.695000   2.170000 ;
      RECT 13.295000   2.100000 15.695000   2.170000 ;
      RECT 13.295000   2.170000 15.765000   2.240000 ;
      RECT 13.295000   2.170000 15.765000   2.240000 ;
      RECT 13.295000   2.240000 15.835000   2.310000 ;
      RECT 13.295000   2.240000 15.835000   2.310000 ;
      RECT 13.295000   2.310000 15.905000   2.380000 ;
      RECT 13.295000   2.310000 15.905000   2.380000 ;
      RECT 13.295000   2.380000 15.975000   2.435000 ;
      RECT 13.295000   2.380000 15.975000   2.435000 ;
      RECT 13.295000   2.435000 16.030000   2.505000 ;
      RECT 13.295000   2.435000 16.030000   2.505000 ;
      RECT 13.295000   2.505000 16.100000   2.575000 ;
      RECT 13.295000   2.505000 16.100000   2.575000 ;
      RECT 13.295000   2.575000 16.170000   2.645000 ;
      RECT 13.295000   2.575000 16.170000   2.645000 ;
      RECT 13.295000   2.645000 16.240000   2.715000 ;
      RECT 13.295000   2.645000 16.240000   2.715000 ;
      RECT 13.295000   2.715000 16.310000   2.785000 ;
      RECT 13.295000   2.715000 16.310000   2.785000 ;
      RECT 13.295000   2.785000 16.380000   2.855000 ;
      RECT 13.295000   2.785000 16.380000   2.855000 ;
      RECT 13.295000   2.855000 16.450000   2.925000 ;
      RECT 13.295000   2.855000 16.450000   2.925000 ;
      RECT 13.295000   2.925000 16.520000   2.995000 ;
      RECT 13.295000   2.925000 16.520000   2.995000 ;
      RECT 13.295000   2.995000 16.590000   3.065000 ;
      RECT 13.295000   2.995000 16.590000   3.065000 ;
      RECT 13.295000   3.065000 16.660000   3.135000 ;
      RECT 13.295000   3.065000 16.660000   3.135000 ;
      RECT 13.295000   3.135000 16.730000   3.205000 ;
      RECT 13.295000   3.135000 16.730000   3.205000 ;
      RECT 13.295000   3.205000 16.800000   3.220000 ;
      RECT 13.295000   3.205000 16.800000   3.220000 ;
      RECT 13.295000   3.220000 16.815000   5.125000 ;
      RECT 13.305000  39.730000 13.855000  39.800000 ;
      RECT 13.320000  39.520000 13.480000  40.370000 ;
      RECT 13.320000  42.530000 29.845000  42.600000 ;
      RECT 13.320000  42.530000 29.845000  42.600000 ;
      RECT 13.365000   5.125000 16.815000   5.195000 ;
      RECT 13.365000   5.125000 16.815000   5.195000 ;
      RECT 13.375000  39.660000 13.925000  39.730000 ;
      RECT 13.390000  42.460000 29.845000  42.530000 ;
      RECT 13.390000  42.460000 29.845000  42.530000 ;
      RECT 13.435000   5.195000 16.815000   5.265000 ;
      RECT 13.435000   5.195000 16.815000   5.265000 ;
      RECT 13.445000  39.590000 13.995000  39.660000 ;
      RECT 13.460000  42.390000 29.845000  42.460000 ;
      RECT 13.460000  42.390000 29.845000  42.460000 ;
      RECT 13.505000   5.265000 16.815000   5.335000 ;
      RECT 13.505000   5.265000 16.815000   5.335000 ;
      RECT 13.515000  39.520000 14.065000  39.590000 ;
      RECT 13.530000  42.320000 29.845000  42.390000 ;
      RECT 13.530000  42.320000 29.845000  42.390000 ;
      RECT 13.575000   5.335000 16.815000   5.405000 ;
      RECT 13.575000   5.335000 16.815000   5.405000 ;
      RECT 13.585000  39.450000 14.135000  39.520000 ;
      RECT 13.600000  42.250000 29.845000  42.320000 ;
      RECT 13.600000  42.250000 29.845000  42.320000 ;
      RECT 13.645000   5.405000 16.815000   5.475000 ;
      RECT 13.645000   5.405000 16.815000   5.475000 ;
      RECT 13.655000  39.380000 14.205000  39.450000 ;
      RECT 13.670000  42.180000 29.845000  42.250000 ;
      RECT 13.670000  42.180000 29.845000  42.250000 ;
      RECT 13.690000  39.345000 15.195000  39.380000 ;
      RECT 13.715000   5.475000 16.815000   5.545000 ;
      RECT 13.715000   5.475000 16.815000   5.545000 ;
      RECT 13.740000  42.110000 29.845000  42.180000 ;
      RECT 13.740000  42.110000 29.845000  42.180000 ;
      RECT 13.760000  39.275000 15.230000  39.345000 ;
      RECT 13.785000   5.545000 16.815000   5.615000 ;
      RECT 13.785000   5.545000 16.815000   5.615000 ;
      RECT 13.810000  42.040000 29.845000  42.110000 ;
      RECT 13.810000  42.040000 29.845000  42.110000 ;
      RECT 13.830000  39.205000 15.300000  39.275000 ;
      RECT 13.855000   5.615000 16.815000   5.685000 ;
      RECT 13.855000   5.615000 16.815000   5.685000 ;
      RECT 13.880000  41.970000 29.845000  42.040000 ;
      RECT 13.880000  41.970000 29.845000  42.040000 ;
      RECT 13.900000  39.135000 15.370000  39.205000 ;
      RECT 13.910000  47.675000 29.985000  48.515000 ;
      RECT 13.925000   5.685000 16.815000   5.755000 ;
      RECT 13.925000   5.685000 16.815000   5.755000 ;
      RECT 13.950000  41.900000 29.845000  41.970000 ;
      RECT 13.950000  41.900000 29.845000  41.970000 ;
      RECT 13.970000  39.065000 15.440000  39.135000 ;
      RECT 13.995000   5.755000 16.815000   5.825000 ;
      RECT 13.995000   5.755000 16.815000   5.825000 ;
      RECT 14.020000  40.600000 29.985000  41.635000 ;
      RECT 14.020000  41.635000 29.985000  44.005000 ;
      RECT 14.020000  41.830000 29.845000  41.900000 ;
      RECT 14.020000  41.830000 29.845000  41.900000 ;
      RECT 14.035000  47.535000 29.845000  47.605000 ;
      RECT 14.035000  47.535000 29.845000  47.605000 ;
      RECT 14.040000  38.995000 15.510000  39.065000 ;
      RECT 14.065000   5.825000 16.815000   5.895000 ;
      RECT 14.065000   5.825000 16.815000   5.895000 ;
      RECT 14.090000  41.760000 29.845000  41.830000 ;
      RECT 14.090000  41.760000 29.845000  41.830000 ;
      RECT 14.105000  47.605000 29.845000  47.675000 ;
      RECT 14.105000  47.605000 29.845000  47.675000 ;
      RECT 14.110000  38.925000 15.580000  38.995000 ;
      RECT 14.135000   5.895000 16.815000   5.965000 ;
      RECT 14.135000   5.895000 16.815000   5.965000 ;
      RECT 14.160000  40.655000 29.845000  41.690000 ;
      RECT 14.160000  41.690000 29.845000  41.760000 ;
      RECT 14.160000  41.690000 29.845000  41.760000 ;
      RECT 14.175000  47.675000 29.845000  47.745000 ;
      RECT 14.175000  47.675000 29.845000  47.745000 ;
      RECT 14.180000  38.855000 15.650000  38.925000 ;
      RECT 14.195000  40.620000 29.845000  40.655000 ;
      RECT 14.195000  40.620000 29.845000  40.655000 ;
      RECT 14.205000   5.965000 16.815000   6.035000 ;
      RECT 14.205000   5.965000 16.815000   6.035000 ;
      RECT 14.245000  47.745000 29.845000  47.815000 ;
      RECT 14.245000  47.745000 29.845000  47.815000 ;
      RECT 14.250000  38.785000 15.720000  38.855000 ;
      RECT 14.265000  40.550000 29.845000  40.620000 ;
      RECT 14.265000  40.550000 29.845000  40.620000 ;
      RECT 14.275000   6.035000 16.815000   6.105000 ;
      RECT 14.275000   6.035000 16.815000   6.105000 ;
      RECT 14.315000  47.815000 29.845000  47.885000 ;
      RECT 14.315000  47.815000 29.845000  47.885000 ;
      RECT 14.320000  38.715000 15.790000  38.785000 ;
      RECT 14.335000  40.480000 29.845000  40.550000 ;
      RECT 14.335000  40.480000 29.845000  40.550000 ;
      RECT 14.345000   6.105000 16.815000   6.175000 ;
      RECT 14.345000   6.105000 16.815000   6.175000 ;
      RECT 14.370000   6.395000 16.955000   6.615000 ;
      RECT 14.370000   6.615000 16.470000   7.100000 ;
      RECT 14.370000   7.100000 16.470000  11.600000 ;
      RECT 14.370000  11.600000 16.565000  11.695000 ;
      RECT 14.370000  11.695000 16.565000  12.320000 ;
      RECT 14.370000  12.320000 16.470000  12.415000 ;
      RECT 14.370000  12.415000 16.470000  18.055000 ;
      RECT 14.370000  18.055000 16.470000  19.470000 ;
      RECT 14.385000  47.885000 29.845000  47.955000 ;
      RECT 14.385000  47.885000 29.845000  47.955000 ;
      RECT 14.390000  38.645000 15.860000  38.715000 ;
      RECT 14.405000  40.410000 29.845000  40.480000 ;
      RECT 14.405000  40.410000 29.845000  40.480000 ;
      RECT 14.415000   6.175000 16.815000   6.245000 ;
      RECT 14.415000   6.175000 16.815000   6.245000 ;
      RECT 14.455000  47.955000 29.845000  48.025000 ;
      RECT 14.455000  47.955000 29.845000  48.025000 ;
      RECT 14.460000  38.575000 15.930000  38.645000 ;
      RECT 14.475000  40.340000 29.845000  40.410000 ;
      RECT 14.475000  40.340000 29.845000  40.410000 ;
      RECT 14.485000   6.245000 16.815000   6.315000 ;
      RECT 14.485000   6.245000 16.815000   6.315000 ;
      RECT 14.510000   6.315000 16.815000   6.340000 ;
      RECT 14.510000   6.315000 16.815000   6.340000 ;
      RECT 14.510000   6.560000 16.745000   6.630000 ;
      RECT 14.510000   6.630000 16.675000   6.700000 ;
      RECT 14.510000   6.700000 16.605000   6.770000 ;
      RECT 14.510000   6.770000 16.535000   6.840000 ;
      RECT 14.510000   6.840000 16.465000   6.910000 ;
      RECT 14.510000   6.910000 16.395000   6.980000 ;
      RECT 14.510000   6.980000 16.330000   7.045000 ;
      RECT 14.510000   7.045000 16.330000  11.655000 ;
      RECT 14.510000  11.655000 16.330000  11.705000 ;
      RECT 14.510000  11.705000 16.380000  11.750000 ;
      RECT 14.510000  11.750000 16.425000  12.265000 ;
      RECT 14.510000  12.265000 16.380000  12.310000 ;
      RECT 14.510000  12.310000 16.335000  12.355000 ;
      RECT 14.510000  12.355000 16.330000  12.360000 ;
      RECT 14.510000  12.360000 16.330000  18.000000 ;
      RECT 14.525000  48.025000 29.845000  48.095000 ;
      RECT 14.525000  48.025000 29.845000  48.095000 ;
      RECT 14.530000  38.505000 16.000000  38.575000 ;
      RECT 14.545000  40.270000 29.845000  40.340000 ;
      RECT 14.545000  40.270000 29.845000  40.340000 ;
      RECT 14.560000  40.060000 29.985000  40.600000 ;
      RECT 14.580000   6.340000 16.815000   6.410000 ;
      RECT 14.580000   6.340000 16.815000   6.410000 ;
      RECT 14.580000  18.000000 16.330000  18.070000 ;
      RECT 14.595000  48.095000 29.845000  48.165000 ;
      RECT 14.595000  48.095000 29.845000  48.165000 ;
      RECT 14.600000  38.435000 16.070000  38.505000 ;
      RECT 14.615000  40.200000 29.845000  40.270000 ;
      RECT 14.615000  40.200000 29.845000  40.270000 ;
      RECT 14.650000   6.410000 16.815000   6.480000 ;
      RECT 14.650000   6.410000 16.815000   6.480000 ;
      RECT 14.650000  18.070000 16.330000  18.140000 ;
      RECT 14.665000  48.165000 29.845000  48.235000 ;
      RECT 14.665000  48.165000 29.845000  48.235000 ;
      RECT 14.670000  38.365000 16.140000  38.435000 ;
      RECT 14.720000   6.480000 16.815000   6.550000 ;
      RECT 14.720000   6.480000 16.815000   6.550000 ;
      RECT 14.720000  18.140000 16.330000  18.210000 ;
      RECT 14.730000   6.550000 16.815000   6.560000 ;
      RECT 14.730000   6.550000 16.815000   6.560000 ;
      RECT 14.735000  48.235000 29.845000  48.305000 ;
      RECT 14.735000  48.235000 29.845000  48.305000 ;
      RECT 14.740000  38.295000 16.210000  38.365000 ;
      RECT 14.750000  48.515000 29.985000  51.370000 ;
      RECT 14.750000  51.370000 29.565000  51.790000 ;
      RECT 14.750000  51.790000 24.535000  53.195000 ;
      RECT 14.750000  53.195000 24.535000  56.895000 ;
      RECT 14.750000  56.895000 24.210000  57.220000 ;
      RECT 14.750000  57.220000 22.940000  57.765000 ;
      RECT 14.750000  57.765000 22.940000  57.780000 ;
      RECT 14.765000  57.780000 76.775000  57.990000 ;
      RECT 14.790000  18.210000 16.330000  18.280000 ;
      RECT 14.800000   6.560000 16.745000   6.630000 ;
      RECT 14.800000   6.560000 16.745000   6.630000 ;
      RECT 14.805000  48.305000 29.845000  48.375000 ;
      RECT 14.805000  48.305000 29.845000  48.375000 ;
      RECT 14.810000  38.225000 16.280000  38.295000 ;
      RECT 14.860000  18.280000 16.330000  18.350000 ;
      RECT 14.870000   6.630000 16.675000   6.700000 ;
      RECT 14.870000   6.630000 16.675000   6.700000 ;
      RECT 14.875000  48.375000 29.845000  48.445000 ;
      RECT 14.875000  48.375000 29.845000  48.445000 ;
      RECT 14.880000  38.155000 16.350000  38.225000 ;
      RECT 14.890000  48.445000 29.845000  48.460000 ;
      RECT 14.890000  48.445000 29.845000  48.460000 ;
      RECT 14.890000  48.460000 29.845000  51.315000 ;
      RECT 14.890000  51.315000 29.775000  51.385000 ;
      RECT 14.890000  51.315000 29.775000  51.385000 ;
      RECT 14.890000  51.385000 29.705000  51.455000 ;
      RECT 14.890000  51.385000 29.705000  51.455000 ;
      RECT 14.890000  51.455000 29.635000  51.525000 ;
      RECT 14.890000  51.455000 29.635000  51.525000 ;
      RECT 14.890000  51.525000 29.565000  51.595000 ;
      RECT 14.890000  51.525000 29.565000  51.595000 ;
      RECT 14.890000  51.595000 29.510000  51.650000 ;
      RECT 14.890000  51.595000 29.510000  51.650000 ;
      RECT 14.890000  51.650000 24.395000  56.840000 ;
      RECT 14.890000  51.650000 25.815000  51.720000 ;
      RECT 14.890000  51.650000 25.815000  51.720000 ;
      RECT 14.890000  51.720000 25.745000  51.790000 ;
      RECT 14.890000  51.720000 25.745000  51.790000 ;
      RECT 14.890000  51.790000 25.675000  51.860000 ;
      RECT 14.890000  51.790000 25.675000  51.860000 ;
      RECT 14.890000  51.860000 25.605000  51.930000 ;
      RECT 14.890000  51.860000 25.605000  51.930000 ;
      RECT 14.890000  51.930000 25.535000  52.000000 ;
      RECT 14.890000  51.930000 25.535000  52.000000 ;
      RECT 14.890000  52.000000 25.465000  52.070000 ;
      RECT 14.890000  52.000000 25.465000  52.070000 ;
      RECT 14.890000  52.070000 25.395000  52.140000 ;
      RECT 14.890000  52.070000 25.395000  52.140000 ;
      RECT 14.890000  52.140000 25.325000  52.210000 ;
      RECT 14.890000  52.140000 25.325000  52.210000 ;
      RECT 14.890000  52.210000 25.255000  52.280000 ;
      RECT 14.890000  52.210000 25.255000  52.280000 ;
      RECT 14.890000  52.280000 25.185000  52.350000 ;
      RECT 14.890000  52.280000 25.185000  52.350000 ;
      RECT 14.890000  52.350000 25.115000  52.420000 ;
      RECT 14.890000  52.350000 25.115000  52.420000 ;
      RECT 14.890000  52.420000 25.045000  52.490000 ;
      RECT 14.890000  52.420000 25.045000  52.490000 ;
      RECT 14.890000  52.490000 24.975000  52.560000 ;
      RECT 14.890000  52.490000 24.975000  52.560000 ;
      RECT 14.890000  52.560000 24.905000  52.630000 ;
      RECT 14.890000  52.560000 24.905000  52.630000 ;
      RECT 14.890000  52.630000 24.835000  52.700000 ;
      RECT 14.890000  52.630000 24.835000  52.700000 ;
      RECT 14.890000  52.700000 24.765000  52.770000 ;
      RECT 14.890000  52.700000 24.765000  52.770000 ;
      RECT 14.890000  52.770000 24.695000  52.840000 ;
      RECT 14.890000  52.770000 24.695000  52.840000 ;
      RECT 14.890000  52.840000 24.625000  52.910000 ;
      RECT 14.890000  52.840000 24.625000  52.910000 ;
      RECT 14.890000  52.910000 24.555000  52.980000 ;
      RECT 14.890000  52.910000 24.555000  52.980000 ;
      RECT 14.890000  52.980000 24.485000  53.050000 ;
      RECT 14.890000  52.980000 24.485000  53.050000 ;
      RECT 14.890000  53.050000 24.415000  53.120000 ;
      RECT 14.890000  53.050000 24.415000  53.120000 ;
      RECT 14.890000  53.120000 24.395000  53.140000 ;
      RECT 14.890000  53.120000 24.395000  53.140000 ;
      RECT 14.890000  53.140000 24.395000  56.840000 ;
      RECT 14.890000  56.840000 24.325000  56.910000 ;
      RECT 14.890000  56.840000 24.325000  56.910000 ;
      RECT 14.890000  56.910000 24.255000  56.980000 ;
      RECT 14.890000  56.910000 24.255000  56.980000 ;
      RECT 14.890000  56.980000 24.185000  57.050000 ;
      RECT 14.890000  56.980000 24.185000  57.050000 ;
      RECT 14.890000  57.050000 24.155000  57.080000 ;
      RECT 14.890000  57.050000 24.155000  57.080000 ;
      RECT 14.890000  57.080000 22.800000  57.710000 ;
      RECT 14.930000  18.350000 16.330000  18.420000 ;
      RECT 14.940000   6.700000 16.605000   6.770000 ;
      RECT 14.940000   6.700000 16.605000   6.770000 ;
      RECT 14.950000  38.085000 16.420000  38.155000 ;
      RECT 14.960000  57.710000 22.800000  57.780000 ;
      RECT 14.960000  57.710000 22.800000  57.780000 ;
      RECT 14.975000  57.990000 76.775000  58.450000 ;
      RECT 15.000000  18.420000 16.330000  18.490000 ;
      RECT 15.010000   6.770000 16.535000   6.840000 ;
      RECT 15.010000   6.770000 16.535000   6.840000 ;
      RECT 15.020000  38.015000 16.490000  38.085000 ;
      RECT 15.030000  57.780000 22.800000  57.850000 ;
      RECT 15.030000  57.780000 22.800000  57.850000 ;
      RECT 15.070000  18.490000 16.330000  18.560000 ;
      RECT 15.080000   6.840000 16.465000   6.910000 ;
      RECT 15.080000   6.840000 16.465000   6.910000 ;
      RECT 15.090000  37.945000 16.560000  38.015000 ;
      RECT 15.100000  57.850000 22.800000  57.920000 ;
      RECT 15.100000  57.850000 22.800000  57.920000 ;
      RECT 15.105000  57.920000 76.635000  57.925000 ;
      RECT 15.105000  57.920000 76.635000  57.925000 ;
      RECT 15.110000  57.925000 76.635000  57.930000 ;
      RECT 15.110000  57.925000 76.635000  57.930000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.920000 76.635000  73.500000 ;
      RECT 15.115000  57.930000 76.635000  57.935000 ;
      RECT 15.115000  57.930000 76.635000  57.935000 ;
      RECT 15.115000  57.935000 76.635000  58.590000 ;
      RECT 15.140000  18.560000 16.330000  18.630000 ;
      RECT 15.150000   6.910000 16.395000   6.980000 ;
      RECT 15.150000   6.910000 16.395000   6.980000 ;
      RECT 15.160000  37.875000 16.630000  37.945000 ;
      RECT 15.210000  18.630000 16.330000  18.700000 ;
      RECT 15.215000   6.980000 16.330000   7.045000 ;
      RECT 15.215000   6.980000 16.330000   7.045000 ;
      RECT 15.230000  37.805000 16.700000  37.875000 ;
      RECT 15.280000  18.700000 16.330000  18.770000 ;
      RECT 15.300000  37.735000 16.770000  37.805000 ;
      RECT 15.350000  18.770000 16.330000  18.840000 ;
      RECT 15.370000  32.130000 16.225000  34.380000 ;
      RECT 15.370000  34.380000 17.435000  35.590000 ;
      RECT 15.370000  35.590000 17.435000  37.335000 ;
      RECT 15.370000  37.335000 17.305000  37.470000 ;
      RECT 15.370000  37.665000 16.840000  37.735000 ;
      RECT 15.420000  18.840000 16.330000  18.910000 ;
      RECT 15.440000  37.595000 16.910000  37.665000 ;
      RECT 15.490000  18.910000 16.330000  18.980000 ;
      RECT 15.510000  32.185000 16.085000  34.435000 ;
      RECT 15.510000  34.435000 16.085000  34.505000 ;
      RECT 15.510000  34.505000 16.155000  34.575000 ;
      RECT 15.510000  34.575000 16.225000  34.645000 ;
      RECT 15.510000  34.645000 16.295000  34.715000 ;
      RECT 15.510000  34.715000 16.365000  34.785000 ;
      RECT 15.510000  34.785000 16.435000  34.855000 ;
      RECT 15.510000  34.855000 16.505000  34.925000 ;
      RECT 15.510000  34.925000 16.575000  34.995000 ;
      RECT 15.510000  34.995000 16.645000  35.065000 ;
      RECT 15.510000  35.065000 16.715000  35.135000 ;
      RECT 15.510000  35.135000 16.785000  35.205000 ;
      RECT 15.510000  35.205000 16.855000  35.275000 ;
      RECT 15.510000  35.275000 16.925000  35.345000 ;
      RECT 15.510000  35.345000 16.995000  35.415000 ;
      RECT 15.510000  35.415000 17.065000  35.485000 ;
      RECT 15.510000  35.485000 17.135000  35.555000 ;
      RECT 15.510000  35.555000 17.205000  35.625000 ;
      RECT 15.510000  35.625000 17.275000  35.645000 ;
      RECT 15.510000  35.645000 17.295000  37.280000 ;
      RECT 15.510000  37.280000 17.225000  37.350000 ;
      RECT 15.510000  37.350000 17.155000  37.420000 ;
      RECT 15.510000  37.420000 17.085000  37.490000 ;
      RECT 15.510000  37.490000 17.050000  37.525000 ;
      RECT 15.510000  37.525000 16.980000  37.595000 ;
      RECT 15.560000  18.980000 16.330000  19.050000 ;
      RECT 15.575000  32.120000 16.085000  32.185000 ;
      RECT 15.590000  40.145000 29.845000  40.200000 ;
      RECT 15.590000  40.145000 29.845000  40.200000 ;
      RECT 15.630000  19.050000 16.330000  19.120000 ;
      RECT 15.645000  32.050000 16.085000  32.120000 ;
      RECT 15.660000  40.075000 29.845000  40.145000 ;
      RECT 15.660000  40.075000 29.845000  40.145000 ;
      RECT 15.700000  19.120000 16.330000  19.190000 ;
      RECT 15.715000  31.980000 16.085000  32.050000 ;
      RECT 15.730000  40.005000 29.845000  40.075000 ;
      RECT 15.730000  40.005000 29.845000  40.075000 ;
      RECT 15.770000  19.190000 16.330000  19.260000 ;
      RECT 15.785000  19.470000 16.470000  31.255000 ;
      RECT 15.785000  31.255000 16.225000  31.500000 ;
      RECT 15.785000  31.500000 16.225000  31.715000 ;
      RECT 15.785000  31.715000 16.225000  32.130000 ;
      RECT 15.785000  31.910000 16.085000  31.980000 ;
      RECT 15.800000  39.935000 29.845000  40.005000 ;
      RECT 15.800000  39.935000 29.845000  40.005000 ;
      RECT 15.840000  19.260000 16.330000  19.330000 ;
      RECT 15.855000  31.840000 16.085000  31.910000 ;
      RECT 15.870000  39.865000 29.845000  39.935000 ;
      RECT 15.870000  39.865000 29.845000  39.935000 ;
      RECT 15.910000  19.330000 16.330000  19.400000 ;
      RECT 15.925000  19.400000 16.330000  19.415000 ;
      RECT 15.925000  19.415000 16.330000  31.200000 ;
      RECT 15.925000  31.200000 16.260000  31.270000 ;
      RECT 15.925000  31.270000 16.190000  31.340000 ;
      RECT 15.925000  31.340000 16.120000  31.410000 ;
      RECT 15.925000  31.410000 16.085000  31.445000 ;
      RECT 15.925000  31.445000 16.085000  31.770000 ;
      RECT 15.925000  31.770000 16.085000  31.840000 ;
      RECT 15.940000  39.795000 29.845000  39.865000 ;
      RECT 15.940000  39.795000 29.845000  39.865000 ;
      RECT 16.010000  39.725000 29.845000  39.795000 ;
      RECT 16.010000  39.725000 29.845000  39.795000 ;
      RECT 16.080000  39.655000 29.845000  39.725000 ;
      RECT 16.080000  39.655000 29.845000  39.725000 ;
      RECT 16.150000  39.585000 29.845000  39.655000 ;
      RECT 16.150000  39.585000 29.845000  39.655000 ;
      RECT 16.220000  39.515000 29.845000  39.585000 ;
      RECT 16.220000  39.515000 29.845000  39.585000 ;
      RECT 16.290000  39.445000 29.845000  39.515000 ;
      RECT 16.290000  39.445000 29.845000  39.515000 ;
      RECT 16.360000  39.375000 29.845000  39.445000 ;
      RECT 16.360000  39.375000 29.845000  39.445000 ;
      RECT 16.430000  39.305000 29.845000  39.375000 ;
      RECT 16.430000  39.305000 29.845000  39.375000 ;
      RECT 16.445000  39.095000 29.985000  40.060000 ;
      RECT 16.500000  39.235000 29.845000  39.305000 ;
      RECT 16.500000  39.235000 29.845000  39.305000 ;
      RECT 16.550000  39.185000 22.815000  39.235000 ;
      RECT 16.550000  39.185000 22.815000  39.235000 ;
      RECT 16.620000  39.115000 22.815000  39.185000 ;
      RECT 16.620000  39.115000 22.815000  39.185000 ;
      RECT 16.690000  39.045000 22.815000  39.115000 ;
      RECT 16.690000  39.045000 22.815000  39.115000 ;
      RECT 16.710000   0.000000 22.215000   2.150000 ;
      RECT 16.710000   2.150000 22.215000   2.935000 ;
      RECT 16.760000  38.975000 22.815000  39.045000 ;
      RECT 16.760000  38.975000 22.815000  39.045000 ;
      RECT 16.765000  31.730000 23.335000  34.150000 ;
      RECT 16.765000  34.150000 23.335000  35.360000 ;
      RECT 16.830000  38.905000 22.815000  38.975000 ;
      RECT 16.830000  38.905000 22.815000  38.975000 ;
      RECT 16.850000   0.000000 22.075000   2.095000 ;
      RECT 16.900000  38.835000 22.815000  38.905000 ;
      RECT 16.900000  38.835000 22.815000  38.905000 ;
      RECT 16.905000  31.785000 23.195000  34.095000 ;
      RECT 16.920000   2.095000 22.075000   2.165000 ;
      RECT 16.920000   2.095000 22.075000   2.165000 ;
      RECT 16.940000  31.750000 23.195000  31.785000 ;
      RECT 16.940000  31.750000 23.195000  31.785000 ;
      RECT 16.970000  38.765000 22.815000  38.835000 ;
      RECT 16.970000  38.765000 22.815000  38.835000 ;
      RECT 16.975000  34.095000 23.195000  34.165000 ;
      RECT 16.975000  34.095000 23.195000  34.165000 ;
      RECT 16.985000  38.555000 22.955000  39.095000 ;
      RECT 16.990000   2.165000 22.075000   2.235000 ;
      RECT 16.990000   2.165000 22.075000   2.235000 ;
      RECT 17.010000   7.330000 22.625000  14.545000 ;
      RECT 17.010000  14.545000 23.515000  15.435000 ;
      RECT 17.010000  15.435000 23.515000  24.940000 ;
      RECT 17.010000  24.940000 23.335000  25.120000 ;
      RECT 17.010000  25.120000 23.335000  31.485000 ;
      RECT 17.010000  31.485000 23.335000  31.730000 ;
      RECT 17.010000  31.680000 23.195000  31.750000 ;
      RECT 17.010000  31.680000 23.195000  31.750000 ;
      RECT 17.040000  38.695000 22.815000  38.765000 ;
      RECT 17.040000  38.695000 22.815000  38.765000 ;
      RECT 17.045000  34.165000 23.195000  34.235000 ;
      RECT 17.045000  34.165000 23.195000  34.235000 ;
      RECT 17.060000   2.235000 22.075000   2.305000 ;
      RECT 17.060000   2.235000 22.075000   2.305000 ;
      RECT 17.080000  31.610000 23.195000  31.680000 ;
      RECT 17.080000  31.610000 23.195000  31.680000 ;
      RECT 17.110000  38.625000 22.815000  38.695000 ;
      RECT 17.110000  38.625000 22.815000  38.695000 ;
      RECT 17.115000  34.235000 23.195000  34.305000 ;
      RECT 17.115000  34.235000 23.195000  34.305000 ;
      RECT 17.130000   2.305000 22.075000   2.375000 ;
      RECT 17.130000   2.305000 22.075000   2.375000 ;
      RECT 17.150000   7.385000 22.485000  14.600000 ;
      RECT 17.150000   7.385000 22.485000  15.490000 ;
      RECT 17.150000  14.600000 22.485000  14.670000 ;
      RECT 17.150000  14.600000 22.485000  14.670000 ;
      RECT 17.150000  14.670000 22.555000  14.740000 ;
      RECT 17.150000  14.670000 22.555000  14.740000 ;
      RECT 17.150000  14.740000 22.625000  14.810000 ;
      RECT 17.150000  14.740000 22.625000  14.810000 ;
      RECT 17.150000  14.810000 22.695000  14.880000 ;
      RECT 17.150000  14.810000 22.695000  14.880000 ;
      RECT 17.150000  14.880000 22.765000  14.950000 ;
      RECT 17.150000  14.880000 22.765000  14.950000 ;
      RECT 17.150000  14.950000 22.835000  15.020000 ;
      RECT 17.150000  14.950000 22.835000  15.020000 ;
      RECT 17.150000  15.020000 22.905000  15.090000 ;
      RECT 17.150000  15.020000 22.905000  15.090000 ;
      RECT 17.150000  15.090000 22.975000  15.160000 ;
      RECT 17.150000  15.090000 22.975000  15.160000 ;
      RECT 17.150000  15.160000 23.045000  15.230000 ;
      RECT 17.150000  15.160000 23.045000  15.230000 ;
      RECT 17.150000  15.230000 23.115000  15.300000 ;
      RECT 17.150000  15.230000 23.115000  15.300000 ;
      RECT 17.150000  15.300000 23.185000  15.370000 ;
      RECT 17.150000  15.300000 23.185000  15.370000 ;
      RECT 17.150000  15.370000 23.255000  15.440000 ;
      RECT 17.150000  15.370000 23.255000  15.440000 ;
      RECT 17.150000  15.440000 23.325000  15.490000 ;
      RECT 17.150000  15.440000 23.325000  15.490000 ;
      RECT 17.150000  15.490000 23.375000  24.885000 ;
      RECT 17.150000  24.885000 23.305000  24.955000 ;
      RECT 17.150000  24.885000 23.305000  24.955000 ;
      RECT 17.150000  24.955000 23.235000  25.025000 ;
      RECT 17.150000  24.955000 23.235000  25.025000 ;
      RECT 17.150000  25.025000 23.195000  25.065000 ;
      RECT 17.150000  25.025000 23.195000  25.065000 ;
      RECT 17.150000  25.065000 23.195000  31.540000 ;
      RECT 17.150000  31.540000 23.195000  31.610000 ;
      RECT 17.150000  31.540000 23.195000  31.610000 ;
      RECT 17.165000   7.370000 22.485000   7.385000 ;
      RECT 17.165000   7.370000 22.485000   7.385000 ;
      RECT 17.180000  38.355000 23.135000  38.555000 ;
      RECT 17.180000  38.555000 22.815000  38.625000 ;
      RECT 17.180000  38.555000 22.815000  38.625000 ;
      RECT 17.185000  34.305000 23.195000  34.375000 ;
      RECT 17.185000  34.305000 23.195000  34.375000 ;
      RECT 17.200000   2.375000 22.075000   2.445000 ;
      RECT 17.200000   2.375000 22.075000   2.445000 ;
      RECT 17.235000   7.300000 22.485000   7.370000 ;
      RECT 17.235000   7.300000 22.485000   7.370000 ;
      RECT 17.250000  38.485000 22.815000  38.555000 ;
      RECT 17.250000  38.485000 22.815000  38.555000 ;
      RECT 17.255000  34.375000 23.195000  34.445000 ;
      RECT 17.255000  34.375000 23.195000  34.445000 ;
      RECT 17.270000   2.445000 22.075000   2.515000 ;
      RECT 17.270000   2.445000 22.075000   2.515000 ;
      RECT 17.305000   7.230000 22.485000   7.300000 ;
      RECT 17.305000   7.230000 22.485000   7.300000 ;
      RECT 17.320000  38.415000 22.815000  38.485000 ;
      RECT 17.320000  38.415000 22.815000  38.485000 ;
      RECT 17.325000  34.445000 23.195000  34.515000 ;
      RECT 17.325000  34.445000 23.195000  34.515000 ;
      RECT 17.340000   2.515000 22.075000   2.585000 ;
      RECT 17.340000   2.515000 22.075000   2.585000 ;
      RECT 17.375000   7.160000 22.485000   7.230000 ;
      RECT 17.375000   7.160000 22.485000   7.230000 ;
      RECT 17.380000  38.355000 23.080000  38.415000 ;
      RECT 17.380000  38.355000 23.080000  38.415000 ;
      RECT 17.395000  34.515000 23.195000  34.585000 ;
      RECT 17.395000  34.515000 23.195000  34.585000 ;
      RECT 17.410000   2.585000 22.075000   2.655000 ;
      RECT 17.410000   2.585000 22.075000   2.655000 ;
      RECT 17.435000  38.300000 23.140000  38.355000 ;
      RECT 17.435000  38.300000 23.140000  38.355000 ;
      RECT 17.445000   6.895000 22.625000   7.330000 ;
      RECT 17.445000   7.090000 22.485000   7.160000 ;
      RECT 17.445000   7.090000 22.485000   7.160000 ;
      RECT 17.465000  34.585000 23.195000  34.655000 ;
      RECT 17.465000  34.585000 23.195000  34.655000 ;
      RECT 17.480000   2.655000 22.075000   2.725000 ;
      RECT 17.480000   2.655000 22.075000   2.725000 ;
      RECT 17.485000  38.250000 23.195000  38.300000 ;
      RECT 17.485000  38.250000 23.195000  38.300000 ;
      RECT 17.495000   2.935000 22.215000   6.480000 ;
      RECT 17.495000   6.480000 22.575000   6.845000 ;
      RECT 17.495000   6.845000 22.625000   6.895000 ;
      RECT 17.515000   7.020000 22.485000   7.090000 ;
      RECT 17.515000   7.020000 22.485000   7.090000 ;
      RECT 17.535000  34.655000 23.195000  34.725000 ;
      RECT 17.535000  34.655000 23.195000  34.725000 ;
      RECT 17.550000   2.725000 22.075000   2.795000 ;
      RECT 17.550000   2.725000 22.075000   2.795000 ;
      RECT 17.555000  38.180000 23.195000  38.250000 ;
      RECT 17.555000  38.180000 23.195000  38.250000 ;
      RECT 17.585000   6.950000 22.485000   7.020000 ;
      RECT 17.585000   6.950000 22.485000   7.020000 ;
      RECT 17.605000  34.725000 23.195000  34.795000 ;
      RECT 17.605000  34.725000 23.195000  34.795000 ;
      RECT 17.610000   6.925000 22.460000   6.950000 ;
      RECT 17.610000   6.925000 22.460000   6.950000 ;
      RECT 17.620000   2.795000 22.075000   2.865000 ;
      RECT 17.620000   2.795000 22.075000   2.865000 ;
      RECT 17.625000  38.110000 23.195000  38.180000 ;
      RECT 17.625000  38.110000 23.195000  38.180000 ;
      RECT 17.635000   0.000000 22.075000   6.540000 ;
      RECT 17.635000   0.000000 22.075000   6.540000 ;
      RECT 17.635000   2.865000 22.075000   2.880000 ;
      RECT 17.635000   2.865000 22.075000   2.880000 ;
      RECT 17.635000   2.880000 22.075000   6.540000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   2.880000 22.075000   6.900000 ;
      RECT 17.635000   6.540000 22.075000   6.610000 ;
      RECT 17.635000   6.540000 22.075000   6.610000 ;
      RECT 17.635000   6.610000 22.145000   6.680000 ;
      RECT 17.635000   6.610000 22.145000   6.680000 ;
      RECT 17.635000   6.680000 22.215000   6.750000 ;
      RECT 17.635000   6.680000 22.215000   6.750000 ;
      RECT 17.635000   6.750000 22.285000   6.820000 ;
      RECT 17.635000   6.750000 22.285000   6.820000 ;
      RECT 17.635000   6.820000 22.355000   6.890000 ;
      RECT 17.635000   6.820000 22.355000   6.890000 ;
      RECT 17.635000   6.890000 22.425000   6.900000 ;
      RECT 17.635000   6.890000 22.425000   6.900000 ;
      RECT 17.635000   6.900000 22.435000   6.925000 ;
      RECT 17.635000   6.900000 22.435000   6.925000 ;
      RECT 17.675000  34.795000 23.195000  34.865000 ;
      RECT 17.675000  34.795000 23.195000  34.865000 ;
      RECT 17.695000  38.040000 23.195000  38.110000 ;
      RECT 17.695000  38.040000 23.195000  38.110000 ;
      RECT 17.745000  34.865000 23.195000  34.935000 ;
      RECT 17.745000  34.865000 23.195000  34.935000 ;
      RECT 17.765000  37.970000 23.195000  38.040000 ;
      RECT 17.765000  37.970000 23.195000  38.040000 ;
      RECT 17.815000  34.935000 23.195000  35.005000 ;
      RECT 17.815000  34.935000 23.195000  35.005000 ;
      RECT 17.835000  37.900000 23.195000  37.970000 ;
      RECT 17.835000  37.900000 23.195000  37.970000 ;
      RECT 17.885000  35.005000 23.195000  35.075000 ;
      RECT 17.885000  35.005000 23.195000  35.075000 ;
      RECT 17.905000  37.830000 23.195000  37.900000 ;
      RECT 17.905000  37.830000 23.195000  37.900000 ;
      RECT 17.955000  35.075000 23.195000  35.145000 ;
      RECT 17.955000  35.075000 23.195000  35.145000 ;
      RECT 17.975000  35.360000 23.335000  37.565000 ;
      RECT 17.975000  37.565000 23.335000  38.355000 ;
      RECT 17.975000  37.760000 23.195000  37.830000 ;
      RECT 17.975000  37.760000 23.195000  37.830000 ;
      RECT 18.025000  35.145000 23.195000  35.215000 ;
      RECT 18.025000  35.145000 23.195000  35.215000 ;
      RECT 18.045000  37.690000 23.195000  37.760000 ;
      RECT 18.045000  37.690000 23.195000  37.760000 ;
      RECT 18.095000  35.215000 23.195000  35.285000 ;
      RECT 18.095000  35.215000 23.195000  35.285000 ;
      RECT 18.115000  31.540000 23.195000  37.620000 ;
      RECT 18.115000  35.285000 23.195000  35.305000 ;
      RECT 18.115000  35.285000 23.195000  35.305000 ;
      RECT 18.115000  35.305000 23.195000  37.620000 ;
      RECT 18.115000  37.620000 23.195000  37.690000 ;
      RECT 18.115000  37.620000 23.195000  37.690000 ;
      RECT 22.755000   0.000000 26.460000   1.835000 ;
      RECT 22.755000   1.835000 28.350000   4.130000 ;
      RECT 22.755000   4.130000 29.070000   4.850000 ;
      RECT 22.755000   4.850000 29.070000   6.255000 ;
      RECT 22.755000   6.255000 29.070000   6.665000 ;
      RECT 22.895000   0.000000 26.320000   1.975000 ;
      RECT 22.895000   0.000000 26.320000   4.185000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   0.000000 26.320000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   4.185000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   1.975000 28.210000   6.200000 ;
      RECT 22.895000   4.185000 28.210000   4.255000 ;
      RECT 22.895000   4.185000 28.210000   4.255000 ;
      RECT 22.895000   4.255000 28.280000   4.325000 ;
      RECT 22.895000   4.255000 28.280000   4.325000 ;
      RECT 22.895000   4.325000 28.350000   4.395000 ;
      RECT 22.895000   4.325000 28.350000   4.395000 ;
      RECT 22.895000   4.395000 28.420000   4.465000 ;
      RECT 22.895000   4.395000 28.420000   4.465000 ;
      RECT 22.895000   4.465000 28.490000   4.535000 ;
      RECT 22.895000   4.465000 28.490000   4.535000 ;
      RECT 22.895000   4.535000 28.560000   4.605000 ;
      RECT 22.895000   4.535000 28.560000   4.605000 ;
      RECT 22.895000   4.605000 28.630000   4.675000 ;
      RECT 22.895000   4.605000 28.630000   4.675000 ;
      RECT 22.895000   4.675000 28.700000   4.745000 ;
      RECT 22.895000   4.675000 28.700000   4.745000 ;
      RECT 22.895000   4.745000 28.770000   4.815000 ;
      RECT 22.895000   4.745000 28.770000   4.815000 ;
      RECT 22.895000   4.815000 28.840000   4.885000 ;
      RECT 22.895000   4.815000 28.840000   4.885000 ;
      RECT 22.895000   4.885000 28.910000   4.905000 ;
      RECT 22.895000   4.885000 28.910000   4.905000 ;
      RECT 22.895000   4.905000 28.930000   6.200000 ;
      RECT 22.965000   6.200000 28.930000   6.270000 ;
      RECT 22.965000   6.200000 28.930000   6.270000 ;
      RECT 23.035000   6.270000 28.930000   6.340000 ;
      RECT 23.035000   6.270000 28.930000   6.340000 ;
      RECT 23.105000   6.340000 28.930000   6.410000 ;
      RECT 23.105000   6.340000 28.930000   6.410000 ;
      RECT 23.165000   6.665000 29.070000   6.920000 ;
      RECT 23.165000   6.920000 31.550000  14.315000 ;
      RECT 23.165000  14.315000 31.550000  15.205000 ;
      RECT 23.175000   6.410000 28.930000   6.480000 ;
      RECT 23.175000   6.410000 28.930000   6.480000 ;
      RECT 23.245000   6.480000 28.930000   6.550000 ;
      RECT 23.245000   6.480000 28.930000   6.550000 ;
      RECT 23.305000   6.550000 28.930000   6.610000 ;
      RECT 23.305000   6.550000 28.930000   6.610000 ;
      RECT 23.305000   6.610000 28.930000   7.060000 ;
      RECT 23.305000   7.060000 31.410000  14.260000 ;
      RECT 23.375000  14.260000 31.410000  14.330000 ;
      RECT 23.375000  14.260000 31.410000  14.330000 ;
      RECT 23.445000  14.330000 31.410000  14.400000 ;
      RECT 23.445000  14.330000 31.410000  14.400000 ;
      RECT 23.515000  14.400000 31.410000  14.470000 ;
      RECT 23.515000  14.400000 31.410000  14.470000 ;
      RECT 23.585000  14.470000 31.410000  14.540000 ;
      RECT 23.585000  14.470000 31.410000  14.540000 ;
      RECT 23.655000  14.540000 31.410000  14.610000 ;
      RECT 23.655000  14.540000 31.410000  14.610000 ;
      RECT 23.725000  14.610000 31.410000  14.680000 ;
      RECT 23.725000  14.610000 31.410000  14.680000 ;
      RECT 23.795000  14.680000 31.410000  14.750000 ;
      RECT 23.795000  14.680000 31.410000  14.750000 ;
      RECT 23.865000  14.750000 31.410000  14.820000 ;
      RECT 23.865000  14.750000 31.410000  14.820000 ;
      RECT 23.875000  25.345000 29.985000  36.515000 ;
      RECT 23.875000  36.515000 30.250000  36.780000 ;
      RECT 23.875000  36.780000 30.250000  37.685000 ;
      RECT 23.875000  37.685000 29.985000  37.950000 ;
      RECT 23.875000  37.950000 29.985000  39.095000 ;
      RECT 23.935000  14.820000 31.410000  14.890000 ;
      RECT 23.935000  14.820000 31.410000  14.890000 ;
      RECT 24.005000  14.890000 31.410000  14.960000 ;
      RECT 24.005000  14.890000 31.410000  14.960000 ;
      RECT 24.015000  25.405000 29.845000  37.630000 ;
      RECT 24.015000  36.570000 29.845000  36.640000 ;
      RECT 24.015000  36.570000 29.845000  36.640000 ;
      RECT 24.015000  36.640000 29.915000  36.710000 ;
      RECT 24.015000  36.640000 29.915000  36.710000 ;
      RECT 24.015000  36.710000 29.985000  36.780000 ;
      RECT 24.015000  36.710000 29.985000  36.780000 ;
      RECT 24.015000  36.780000 30.055000  36.835000 ;
      RECT 24.015000  36.780000 30.055000  36.835000 ;
      RECT 24.015000  36.835000 30.110000  37.245000 ;
      RECT 24.015000  37.245000 30.110000  37.630000 ;
      RECT 24.015000  37.630000 30.040000  37.700000 ;
      RECT 24.015000  37.630000 30.040000  37.700000 ;
      RECT 24.015000  37.700000 29.970000  37.770000 ;
      RECT 24.015000  37.700000 29.970000  37.770000 ;
      RECT 24.015000  37.770000 29.900000  37.840000 ;
      RECT 24.015000  37.770000 29.900000  37.840000 ;
      RECT 24.015000  37.840000 29.845000  37.895000 ;
      RECT 24.015000  37.840000 29.845000  37.895000 ;
      RECT 24.015000  37.895000 29.845000  39.235000 ;
      RECT 24.055000  15.205000 31.550000  16.005000 ;
      RECT 24.055000  16.005000 29.985000  17.570000 ;
      RECT 24.055000  17.570000 29.985000  25.165000 ;
      RECT 24.055000  25.165000 29.985000  25.345000 ;
      RECT 24.055000  25.365000 29.845000  25.405000 ;
      RECT 24.055000  25.365000 29.845000  25.405000 ;
      RECT 24.075000  14.960000 31.410000  15.030000 ;
      RECT 24.075000  14.960000 31.410000  15.030000 ;
      RECT 24.125000  25.295000 29.845000  25.365000 ;
      RECT 24.125000  25.295000 29.845000  25.365000 ;
      RECT 24.145000  15.030000 31.410000  15.100000 ;
      RECT 24.145000  15.030000 31.410000  15.100000 ;
      RECT 24.195000  15.100000 31.410000  15.150000 ;
      RECT 24.195000  15.100000 31.410000  15.150000 ;
      RECT 24.195000  15.150000 31.410000  15.950000 ;
      RECT 24.195000  15.950000 29.845000  25.225000 ;
      RECT 24.195000  15.950000 31.340000  16.020000 ;
      RECT 24.195000  15.950000 31.340000  16.020000 ;
      RECT 24.195000  16.020000 31.270000  16.090000 ;
      RECT 24.195000  16.020000 31.270000  16.090000 ;
      RECT 24.195000  16.090000 31.200000  16.160000 ;
      RECT 24.195000  16.090000 31.200000  16.160000 ;
      RECT 24.195000  16.160000 31.130000  16.230000 ;
      RECT 24.195000  16.160000 31.130000  16.230000 ;
      RECT 24.195000  16.230000 31.060000  16.300000 ;
      RECT 24.195000  16.230000 31.060000  16.300000 ;
      RECT 24.195000  16.300000 30.990000  16.370000 ;
      RECT 24.195000  16.300000 30.990000  16.370000 ;
      RECT 24.195000  16.370000 30.920000  16.440000 ;
      RECT 24.195000  16.370000 30.920000  16.440000 ;
      RECT 24.195000  16.440000 30.850000  16.510000 ;
      RECT 24.195000  16.440000 30.850000  16.510000 ;
      RECT 24.195000  16.510000 30.780000  16.580000 ;
      RECT 24.195000  16.510000 30.780000  16.580000 ;
      RECT 24.195000  16.580000 30.710000  16.650000 ;
      RECT 24.195000  16.580000 30.710000  16.650000 ;
      RECT 24.195000  16.650000 30.640000  16.720000 ;
      RECT 24.195000  16.650000 30.640000  16.720000 ;
      RECT 24.195000  16.720000 30.570000  16.790000 ;
      RECT 24.195000  16.720000 30.570000  16.790000 ;
      RECT 24.195000  16.790000 30.500000  16.860000 ;
      RECT 24.195000  16.790000 30.500000  16.860000 ;
      RECT 24.195000  16.860000 30.430000  16.930000 ;
      RECT 24.195000  16.860000 30.430000  16.930000 ;
      RECT 24.195000  16.930000 30.360000  17.000000 ;
      RECT 24.195000  16.930000 30.360000  17.000000 ;
      RECT 24.195000  17.000000 30.290000  17.070000 ;
      RECT 24.195000  17.000000 30.290000  17.070000 ;
      RECT 24.195000  17.070000 30.220000  17.140000 ;
      RECT 24.195000  17.070000 30.220000  17.140000 ;
      RECT 24.195000  17.140000 30.150000  17.210000 ;
      RECT 24.195000  17.140000 30.150000  17.210000 ;
      RECT 24.195000  17.210000 30.080000  17.280000 ;
      RECT 24.195000  17.210000 30.080000  17.280000 ;
      RECT 24.195000  17.280000 30.010000  17.350000 ;
      RECT 24.195000  17.280000 30.010000  17.350000 ;
      RECT 24.195000  17.350000 29.940000  17.420000 ;
      RECT 24.195000  17.350000 29.940000  17.420000 ;
      RECT 24.195000  17.420000 29.870000  17.490000 ;
      RECT 24.195000  17.420000 29.870000  17.490000 ;
      RECT 24.195000  17.490000 29.845000  17.515000 ;
      RECT 24.195000  17.490000 29.845000  17.515000 ;
      RECT 24.195000  17.515000 29.845000  25.225000 ;
      RECT 24.195000  25.225000 29.845000  25.295000 ;
      RECT 24.195000  25.225000 29.845000  25.295000 ;
      RECT 24.535000  57.880000 76.635000  57.920000 ;
      RECT 24.535000  57.880000 76.635000  57.920000 ;
      RECT 24.605000  57.810000 76.635000  57.880000 ;
      RECT 24.605000  57.810000 76.635000  57.880000 ;
      RECT 24.675000  57.740000 76.635000  57.810000 ;
      RECT 24.675000  57.740000 76.635000  57.810000 ;
      RECT 24.745000  57.670000 76.635000  57.740000 ;
      RECT 24.745000  57.670000 76.635000  57.740000 ;
      RECT 24.815000  57.600000 76.635000  57.670000 ;
      RECT 24.815000  57.600000 76.635000  57.670000 ;
      RECT 24.885000  57.530000 76.635000  57.600000 ;
      RECT 24.885000  57.530000 76.635000  57.600000 ;
      RECT 24.955000  57.460000 76.635000  57.530000 ;
      RECT 24.955000  57.460000 76.635000  57.530000 ;
      RECT 25.025000  57.390000 76.635000  57.460000 ;
      RECT 25.025000  57.390000 76.635000  57.460000 ;
      RECT 25.095000  53.425000 76.775000  57.125000 ;
      RECT 25.095000  57.125000 76.775000  57.780000 ;
      RECT 25.095000  57.320000 76.635000  57.390000 ;
      RECT 25.095000  57.320000 76.635000  57.390000 ;
      RECT 25.165000  57.250000 76.635000  57.320000 ;
      RECT 25.165000  57.250000 76.635000  57.320000 ;
      RECT 25.235000  53.480000 76.635000  57.180000 ;
      RECT 25.235000  53.480000 76.635000  57.920000 ;
      RECT 25.235000  53.480000 76.635000  73.500000 ;
      RECT 25.235000  57.180000 76.635000  57.250000 ;
      RECT 25.235000  57.180000 76.635000  57.250000 ;
      RECT 25.260000  53.260000 76.775000  53.425000 ;
      RECT 25.260000  53.455000 76.635000  53.480000 ;
      RECT 25.260000  53.455000 76.635000  53.480000 ;
      RECT 25.330000  53.385000 76.635000  53.455000 ;
      RECT 25.330000  53.385000 76.635000  53.455000 ;
      RECT 25.400000  53.315000 76.635000  53.385000 ;
      RECT 25.400000  53.315000 76.635000  53.385000 ;
      RECT 25.455000  53.260000 76.580000  53.315000 ;
      RECT 25.455000  53.260000 76.580000  53.315000 ;
      RECT 25.525000  53.190000 76.510000  53.260000 ;
      RECT 25.525000  53.190000 76.510000  53.260000 ;
      RECT 25.595000  53.120000 76.440000  53.190000 ;
      RECT 25.595000  53.120000 76.440000  53.190000 ;
      RECT 25.665000  53.050000 76.370000  53.120000 ;
      RECT 25.665000  53.050000 76.370000  53.120000 ;
      RECT 25.735000  52.980000 76.300000  53.050000 ;
      RECT 25.735000  52.980000 76.300000  53.050000 ;
      RECT 25.805000  52.910000 76.230000  52.980000 ;
      RECT 25.805000  52.910000 76.230000  52.980000 ;
      RECT 25.875000  52.840000 76.160000  52.910000 ;
      RECT 25.875000  52.840000 76.160000  52.910000 ;
      RECT 25.945000  52.575000 76.775000  53.260000 ;
      RECT 25.945000  52.770000 76.090000  52.840000 ;
      RECT 25.945000  52.770000 76.090000  52.840000 ;
      RECT 26.015000  52.700000 76.020000  52.770000 ;
      RECT 26.015000  52.700000 76.020000  52.770000 ;
      RECT 26.085000  52.630000 75.950000  52.700000 ;
      RECT 26.085000  52.630000 75.950000  52.700000 ;
      RECT 26.155000  52.560000 75.950000  52.630000 ;
      RECT 26.155000  52.560000 75.950000  52.630000 ;
      RECT 26.165000  52.350000 76.090000  52.575000 ;
      RECT 26.225000  52.490000 75.950000  52.560000 ;
      RECT 26.225000  52.490000 75.950000  52.560000 ;
      RECT 27.000000   0.000000 28.350000   1.835000 ;
      RECT 27.140000   0.000000 28.210000   1.975000 ;
      RECT 28.890000   0.000000 30.610000   2.320000 ;
      RECT 28.890000   2.320000 31.165000   2.880000 ;
      RECT 28.890000   2.880000 31.165000   3.900000 ;
      RECT 28.890000   3.900000 31.165000   4.505000 ;
      RECT 29.030000   0.000000 30.470000   2.380000 ;
      RECT 29.030000   2.380000 30.470000   2.450000 ;
      RECT 29.030000   2.450000 30.540000   2.520000 ;
      RECT 29.030000   2.520000 30.610000   2.590000 ;
      RECT 29.030000   2.590000 30.680000   2.660000 ;
      RECT 29.030000   2.660000 30.750000   2.730000 ;
      RECT 29.030000   2.730000 30.820000   2.800000 ;
      RECT 29.030000   2.800000 30.890000   2.870000 ;
      RECT 29.030000   2.870000 30.960000   2.935000 ;
      RECT 29.030000   2.935000 31.025000   3.845000 ;
      RECT 29.100000   3.845000 31.025000   3.915000 ;
      RECT 29.170000   3.915000 31.025000   3.985000 ;
      RECT 29.240000   3.985000 31.025000   4.055000 ;
      RECT 29.310000   4.055000 31.025000   4.125000 ;
      RECT 29.380000   4.125000 31.025000   4.195000 ;
      RECT 29.450000   4.195000 31.025000   4.265000 ;
      RECT 29.490000   4.505000 31.285000   4.620000 ;
      RECT 29.520000   4.265000 31.025000   4.335000 ;
      RECT 29.590000   4.335000 31.025000   4.405000 ;
      RECT 29.610000   4.620000 31.550000   4.890000 ;
      RECT 29.610000   4.890000 31.550000   6.920000 ;
      RECT 29.660000   4.405000 31.025000   4.475000 ;
      RECT 29.730000   4.475000 31.025000   4.545000 ;
      RECT 29.745000   4.545000 31.025000   4.560000 ;
      RECT 29.750000   4.560000 31.025000   4.565000 ;
      RECT 29.750000   4.565000 31.025000   4.635000 ;
      RECT 29.750000   4.635000 31.100000   4.705000 ;
      RECT 29.750000   4.705000 31.170000   4.775000 ;
      RECT 29.750000   4.775000 31.240000   4.845000 ;
      RECT 29.750000   4.845000 31.310000   4.915000 ;
      RECT 29.750000   4.915000 31.380000   4.945000 ;
      RECT 29.750000   4.945000 31.410000   7.060000 ;
      RECT 29.895000  52.445000 75.950000  52.490000 ;
      RECT 29.895000  52.445000 75.950000  52.490000 ;
      RECT 29.965000  52.375000 75.950000  52.445000 ;
      RECT 29.965000  52.375000 75.950000  52.445000 ;
      RECT 30.035000  52.305000 75.950000  52.375000 ;
      RECT 30.035000  52.305000 75.950000  52.375000 ;
      RECT 30.105000  52.235000 75.950000  52.305000 ;
      RECT 30.105000  52.235000 75.950000  52.305000 ;
      RECT 30.175000  52.165000 75.950000  52.235000 ;
      RECT 30.175000  52.165000 75.950000  52.235000 ;
      RECT 30.245000  52.095000 75.950000  52.165000 ;
      RECT 30.245000  52.095000 75.950000  52.165000 ;
      RECT 30.315000  52.025000 75.950000  52.095000 ;
      RECT 30.315000  52.025000 75.950000  52.095000 ;
      RECT 30.385000  51.955000 75.950000  52.025000 ;
      RECT 30.385000  51.955000 75.950000  52.025000 ;
      RECT 30.455000  51.885000 75.950000  51.955000 ;
      RECT 30.455000  51.885000 75.950000  51.955000 ;
      RECT 30.525000  17.795000 79.180000  36.285000 ;
      RECT 30.525000  36.285000 79.180000  36.550000 ;
      RECT 30.525000  38.180000 79.180000  47.610000 ;
      RECT 30.525000  47.610000 76.090000  50.700000 ;
      RECT 30.525000  50.700000 76.090000  51.620000 ;
      RECT 30.525000  51.620000 76.090000  52.350000 ;
      RECT 30.525000  51.815000 75.950000  51.885000 ;
      RECT 30.525000  51.815000 75.950000  51.885000 ;
      RECT 30.595000  51.745000 75.950000  51.815000 ;
      RECT 30.595000  51.745000 75.950000  51.815000 ;
      RECT 30.665000  17.855000 79.175000  36.230000 ;
      RECT 30.665000  38.235000 79.175000  42.955000 ;
      RECT 30.665000  42.955000 75.950000  52.490000 ;
      RECT 30.665000  42.955000 79.040000  47.555000 ;
      RECT 30.665000  47.555000 75.950000  52.490000 ;
      RECT 30.665000  47.555000 78.970000  47.625000 ;
      RECT 30.665000  47.555000 78.970000  47.625000 ;
      RECT 30.665000  47.625000 78.900000  47.695000 ;
      RECT 30.665000  47.625000 78.900000  47.695000 ;
      RECT 30.665000  47.695000 78.830000  47.765000 ;
      RECT 30.665000  47.695000 78.830000  47.765000 ;
      RECT 30.665000  47.765000 78.760000  47.835000 ;
      RECT 30.665000  47.765000 78.760000  47.835000 ;
      RECT 30.665000  47.835000 78.690000  47.905000 ;
      RECT 30.665000  47.835000 78.690000  47.905000 ;
      RECT 30.665000  47.905000 78.620000  47.975000 ;
      RECT 30.665000  47.905000 78.620000  47.975000 ;
      RECT 30.665000  47.975000 78.550000  48.045000 ;
      RECT 30.665000  47.975000 78.550000  48.045000 ;
      RECT 30.665000  48.045000 78.480000  48.115000 ;
      RECT 30.665000  48.045000 78.480000  48.115000 ;
      RECT 30.665000  48.115000 78.410000  48.185000 ;
      RECT 30.665000  48.115000 78.410000  48.185000 ;
      RECT 30.665000  48.185000 78.340000  48.255000 ;
      RECT 30.665000  48.185000 78.340000  48.255000 ;
      RECT 30.665000  48.255000 78.270000  48.325000 ;
      RECT 30.665000  48.255000 78.270000  48.325000 ;
      RECT 30.665000  48.325000 78.200000  48.395000 ;
      RECT 30.665000  48.325000 78.200000  48.395000 ;
      RECT 30.665000  48.395000 78.130000  48.465000 ;
      RECT 30.665000  48.395000 78.130000  48.465000 ;
      RECT 30.665000  48.465000 78.060000  48.535000 ;
      RECT 30.665000  48.465000 78.060000  48.535000 ;
      RECT 30.665000  48.535000 77.990000  48.605000 ;
      RECT 30.665000  48.535000 77.990000  48.605000 ;
      RECT 30.665000  48.605000 77.920000  48.675000 ;
      RECT 30.665000  48.605000 77.920000  48.675000 ;
      RECT 30.665000  48.675000 77.850000  48.745000 ;
      RECT 30.665000  48.675000 77.850000  48.745000 ;
      RECT 30.665000  48.745000 77.780000  48.815000 ;
      RECT 30.665000  48.745000 77.780000  48.815000 ;
      RECT 30.665000  48.815000 77.710000  48.885000 ;
      RECT 30.665000  48.815000 77.710000  48.885000 ;
      RECT 30.665000  48.885000 77.640000  48.955000 ;
      RECT 30.665000  48.885000 77.640000  48.955000 ;
      RECT 30.665000  48.955000 77.570000  49.025000 ;
      RECT 30.665000  48.955000 77.570000  49.025000 ;
      RECT 30.665000  49.025000 77.500000  49.095000 ;
      RECT 30.665000  49.025000 77.500000  49.095000 ;
      RECT 30.665000  49.095000 77.430000  49.165000 ;
      RECT 30.665000  49.095000 77.430000  49.165000 ;
      RECT 30.665000  49.165000 77.360000  49.235000 ;
      RECT 30.665000  49.165000 77.360000  49.235000 ;
      RECT 30.665000  49.235000 77.290000  49.305000 ;
      RECT 30.665000  49.235000 77.290000  49.305000 ;
      RECT 30.665000  49.305000 77.220000  49.375000 ;
      RECT 30.665000  49.305000 77.220000  49.375000 ;
      RECT 30.665000  49.375000 77.150000  49.445000 ;
      RECT 30.665000  49.375000 77.150000  49.445000 ;
      RECT 30.665000  49.445000 77.080000  49.515000 ;
      RECT 30.665000  49.445000 77.080000  49.515000 ;
      RECT 30.665000  49.515000 77.010000  49.585000 ;
      RECT 30.665000  49.515000 77.010000  49.585000 ;
      RECT 30.665000  49.585000 76.940000  49.655000 ;
      RECT 30.665000  49.585000 76.940000  49.655000 ;
      RECT 30.665000  49.655000 76.870000  49.725000 ;
      RECT 30.665000  49.655000 76.870000  49.725000 ;
      RECT 30.665000  49.725000 76.800000  49.795000 ;
      RECT 30.665000  49.725000 76.800000  49.795000 ;
      RECT 30.665000  49.795000 76.730000  49.865000 ;
      RECT 30.665000  49.795000 76.730000  49.865000 ;
      RECT 30.665000  49.865000 76.660000  49.935000 ;
      RECT 30.665000  49.865000 76.660000  49.935000 ;
      RECT 30.665000  49.935000 76.590000  50.005000 ;
      RECT 30.665000  49.935000 76.590000  50.005000 ;
      RECT 30.665000  50.005000 76.520000  50.075000 ;
      RECT 30.665000  50.005000 76.520000  50.075000 ;
      RECT 30.665000  50.075000 76.450000  50.145000 ;
      RECT 30.665000  50.075000 76.450000  50.145000 ;
      RECT 30.665000  50.145000 76.380000  50.215000 ;
      RECT 30.665000  50.145000 76.380000  50.215000 ;
      RECT 30.665000  50.215000 76.310000  50.285000 ;
      RECT 30.665000  50.215000 76.310000  50.285000 ;
      RECT 30.665000  50.285000 76.240000  50.355000 ;
      RECT 30.665000  50.285000 76.240000  50.355000 ;
      RECT 30.665000  50.355000 76.170000  50.425000 ;
      RECT 30.665000  50.355000 76.170000  50.425000 ;
      RECT 30.665000  50.425000 76.100000  50.495000 ;
      RECT 30.665000  50.425000 76.100000  50.495000 ;
      RECT 30.665000  50.495000 76.030000  50.565000 ;
      RECT 30.665000  50.495000 76.030000  50.565000 ;
      RECT 30.665000  50.565000 75.960000  50.635000 ;
      RECT 30.665000  50.565000 75.960000  50.635000 ;
      RECT 30.665000  50.635000 75.950000  50.645000 ;
      RECT 30.665000  50.635000 75.950000  50.645000 ;
      RECT 30.665000  50.645000 75.950000  51.675000 ;
      RECT 30.665000  51.675000 75.950000  51.745000 ;
      RECT 30.665000  51.675000 75.950000  51.745000 ;
      RECT 30.715000  17.805000 79.175000  17.855000 ;
      RECT 30.715000  17.805000 79.175000  17.855000 ;
      RECT 30.720000  38.180000 79.175000  38.235000 ;
      RECT 30.720000  38.180000 79.175000  38.235000 ;
      RECT 30.735000  36.230000 79.175000  36.300000 ;
      RECT 30.735000  36.230000 79.175000  36.300000 ;
      RECT 30.785000  17.735000 79.175000  17.805000 ;
      RECT 30.785000  17.735000 79.175000  17.805000 ;
      RECT 30.790000  36.550000 79.180000  37.915000 ;
      RECT 30.790000  37.915000 79.180000  38.180000 ;
      RECT 30.790000  38.110000 79.175000  38.180000 ;
      RECT 30.790000  38.110000 79.175000  38.180000 ;
      RECT 30.805000  36.300000 79.175000  36.370000 ;
      RECT 30.805000  36.300000 79.175000  36.370000 ;
      RECT 30.855000  17.665000 79.175000  17.735000 ;
      RECT 30.855000  17.665000 79.175000  17.735000 ;
      RECT 30.860000  38.040000 79.175000  38.110000 ;
      RECT 30.860000  38.040000 79.175000  38.110000 ;
      RECT 30.875000  36.370000 79.175000  36.440000 ;
      RECT 30.875000  36.370000 79.175000  36.440000 ;
      RECT 30.925000  17.595000 79.175000  17.665000 ;
      RECT 30.925000  17.595000 79.175000  17.665000 ;
      RECT 30.930000  17.855000 79.175000  42.955000 ;
      RECT 30.930000  36.440000 79.175000  36.495000 ;
      RECT 30.930000  36.440000 79.175000  36.495000 ;
      RECT 30.930000  37.970000 79.175000  38.040000 ;
      RECT 30.930000  37.970000 79.175000  38.040000 ;
      RECT 30.995000  17.525000 79.175000  17.595000 ;
      RECT 30.995000  17.525000 79.175000  17.595000 ;
      RECT 31.065000  17.455000 79.175000  17.525000 ;
      RECT 31.065000  17.455000 79.175000  17.525000 ;
      RECT 31.135000  17.385000 79.175000  17.455000 ;
      RECT 31.135000  17.385000 79.175000  17.455000 ;
      RECT 31.150000   0.000000 31.675000   2.095000 ;
      RECT 31.150000   2.095000 31.675000   2.620000 ;
      RECT 31.205000  17.315000 79.175000  17.385000 ;
      RECT 31.205000  17.315000 79.175000  17.385000 ;
      RECT 31.210000  17.310000 79.170000  17.315000 ;
      RECT 31.210000  17.310000 79.170000  17.315000 ;
      RECT 31.235000  17.090000 79.180000  17.795000 ;
      RECT 31.275000  17.245000 79.105000  17.310000 ;
      RECT 31.275000  17.245000 79.105000  17.310000 ;
      RECT 31.290000   0.000000 31.535000   2.040000 ;
      RECT 31.340000  17.180000 79.040000  17.245000 ;
      RECT 31.340000  17.180000 79.040000  17.245000 ;
      RECT 31.355000  17.165000 79.040000  17.180000 ;
      RECT 31.355000  17.165000 79.040000  17.180000 ;
      RECT 31.360000   2.040000 31.535000   2.110000 ;
      RECT 31.375000  17.145000 79.040000  17.165000 ;
      RECT 31.375000  17.145000 79.040000  17.165000 ;
      RECT 31.430000   2.110000 31.535000   2.180000 ;
      RECT 31.435000  17.085000 78.980000  17.145000 ;
      RECT 31.435000  17.085000 78.980000  17.145000 ;
      RECT 31.500000   2.180000 31.535000   2.250000 ;
      RECT 31.505000  17.015000 78.910000  17.085000 ;
      RECT 31.505000  17.015000 78.910000  17.085000 ;
      RECT 31.575000  16.945000 78.840000  17.015000 ;
      RECT 31.575000  16.945000 78.840000  17.015000 ;
      RECT 31.645000  16.875000 78.770000  16.945000 ;
      RECT 31.645000  16.875000 78.770000  16.945000 ;
      RECT 31.705000   4.105000 45.105000   4.275000 ;
      RECT 31.705000   4.275000 45.105000   4.660000 ;
      RECT 31.715000  16.805000 78.700000  16.875000 ;
      RECT 31.715000  16.805000 78.700000  16.875000 ;
      RECT 31.785000  16.735000 78.630000  16.805000 ;
      RECT 31.785000  16.735000 78.630000  16.805000 ;
      RECT 31.855000  16.665000 78.560000  16.735000 ;
      RECT 31.855000  16.665000 78.560000  16.735000 ;
      RECT 31.925000  16.595000 78.490000  16.665000 ;
      RECT 31.925000  16.595000 78.490000  16.665000 ;
      RECT 31.940000   4.245000 44.965000   4.315000 ;
      RECT 31.940000  16.380000 79.180000  17.090000 ;
      RECT 31.995000  16.525000 78.420000  16.595000 ;
      RECT 31.995000  16.525000 78.420000  16.595000 ;
      RECT 32.010000   4.315000 44.965000   4.385000 ;
      RECT 32.020000  16.500000 78.420000  16.525000 ;
      RECT 32.020000  16.500000 78.420000  16.525000 ;
      RECT 32.080000   4.385000 44.965000   4.455000 ;
      RECT 32.090000   4.660000 45.105000   5.145000 ;
      RECT 32.090000   5.145000 45.715000   5.760000 ;
      RECT 32.090000   5.760000 45.715000   6.920000 ;
      RECT 32.090000   6.920000 78.570000  10.110000 ;
      RECT 32.090000  10.110000 78.475000  10.205000 ;
      RECT 32.090000  10.205000 78.475000  16.235000 ;
      RECT 32.090000  16.235000 78.475000  16.380000 ;
      RECT 32.090000  16.430000 78.420000  16.500000 ;
      RECT 32.090000  16.430000 78.420000  16.500000 ;
      RECT 32.150000   4.455000 44.965000   4.525000 ;
      RECT 32.160000  16.360000 78.420000  16.430000 ;
      RECT 32.160000  16.360000 78.420000  16.430000 ;
      RECT 32.215000   0.000000 35.320000   1.840000 ;
      RECT 32.215000   1.840000 34.995000   2.165000 ;
      RECT 32.215000   2.165000 34.995000   4.025000 ;
      RECT 32.215000   4.025000 45.105000   4.105000 ;
      RECT 32.220000   4.525000 44.965000   4.595000 ;
      RECT 32.230000   4.245000 44.965000   4.605000 ;
      RECT 32.230000   4.595000 44.965000   4.605000 ;
      RECT 32.230000   4.605000 44.965000   5.205000 ;
      RECT 32.230000   5.205000 44.965000   5.275000 ;
      RECT 32.230000   5.205000 44.965000   5.275000 ;
      RECT 32.230000   5.275000 45.035000   5.345000 ;
      RECT 32.230000   5.275000 45.035000   5.345000 ;
      RECT 32.230000   5.345000 45.105000   5.415000 ;
      RECT 32.230000   5.345000 45.105000   5.415000 ;
      RECT 32.230000   5.415000 45.175000   5.485000 ;
      RECT 32.230000   5.415000 45.175000   5.485000 ;
      RECT 32.230000   5.485000 45.245000   5.555000 ;
      RECT 32.230000   5.485000 45.245000   5.555000 ;
      RECT 32.230000   5.555000 45.315000   5.625000 ;
      RECT 32.230000   5.555000 45.315000   5.625000 ;
      RECT 32.230000   5.625000 45.385000   5.695000 ;
      RECT 32.230000   5.625000 45.385000   5.695000 ;
      RECT 32.230000   5.695000 45.455000   5.765000 ;
      RECT 32.230000   5.695000 45.455000   5.765000 ;
      RECT 32.230000   5.765000 45.525000   5.815000 ;
      RECT 32.230000   5.765000 45.525000   5.815000 ;
      RECT 32.230000   5.815000 45.575000   7.060000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.420000  16.290000 ;
      RECT 32.230000   7.060000 78.430000   8.230000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.230000 78.430000   8.295000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.295000 78.495000   8.360000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.360000 78.560000   8.365000 ;
      RECT 32.230000   8.365000 78.565000   9.910000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.910000 78.500000   9.975000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000   9.975000 78.435000  10.040000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.040000 78.430000  10.045000 ;
      RECT 32.230000  10.045000 78.430000  10.055000 ;
      RECT 32.230000  10.055000 78.425000  10.060000 ;
      RECT 32.230000  10.055000 78.425000  10.060000 ;
      RECT 32.230000  10.060000 78.420000  10.065000 ;
      RECT 32.230000  10.060000 78.420000  10.065000 ;
      RECT 32.230000  10.065000 78.420000  16.290000 ;
      RECT 32.230000  10.065000 78.420000  17.855000 ;
      RECT 32.230000  16.290000 78.420000  16.360000 ;
      RECT 32.230000  16.290000 78.420000  16.360000 ;
      RECT 32.355000   0.000000 35.180000   1.785000 ;
      RECT 32.355000   1.785000 35.110000   1.855000 ;
      RECT 32.355000   1.855000 35.040000   1.925000 ;
      RECT 32.355000   1.925000 34.970000   1.995000 ;
      RECT 32.355000   1.995000 34.900000   2.065000 ;
      RECT 32.355000   2.065000 34.855000   2.110000 ;
      RECT 32.355000   2.110000 34.855000   4.165000 ;
      RECT 32.355000   4.165000 44.965000   4.245000 ;
      RECT 35.535000   2.390000 38.250000   3.855000 ;
      RECT 35.535000   3.855000 45.105000   4.025000 ;
      RECT 35.675000   2.450000 38.110000   3.995000 ;
      RECT 35.675000   3.995000 44.965000   4.165000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.675000   3.995000 44.965000   7.060000 ;
      RECT 35.720000   2.405000 38.110000   2.450000 ;
      RECT 35.790000   2.335000 38.110000   2.405000 ;
      RECT 35.860000   0.000000 38.250000   2.070000 ;
      RECT 35.860000   2.070000 38.250000   2.390000 ;
      RECT 35.860000   2.265000 38.110000   2.335000 ;
      RECT 35.930000   2.195000 38.110000   2.265000 ;
      RECT 36.000000   0.000000 38.110000   2.125000 ;
      RECT 36.000000   2.125000 38.110000   2.195000 ;
      RECT 38.790000   0.000000 45.105000   3.855000 ;
      RECT 38.930000   0.000000 44.965000   3.995000 ;
      RECT 38.930000   0.000000 44.965000   4.605000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   5.205000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 38.930000   0.000000 44.965000   7.060000 ;
      RECT 45.645000   0.000000 49.715000   0.220000 ;
      RECT 45.645000   0.220000 49.450000   0.485000 ;
      RECT 45.645000   0.485000 49.450000   0.965000 ;
      RECT 45.645000   0.965000 66.400000   1.135000 ;
      RECT 45.645000   1.135000 66.400000   1.615000 ;
      RECT 45.645000   1.615000 68.135000   4.100000 ;
      RECT 45.645000   4.100000 77.010000   4.920000 ;
      RECT 45.645000   4.920000 77.010000   5.375000 ;
      RECT 45.785000   0.000000 49.310000   0.165000 ;
      RECT 45.785000   0.165000 49.310000   0.430000 ;
      RECT 45.785000   0.165000 49.505000   0.235000 ;
      RECT 45.785000   0.235000 49.435000   0.305000 ;
      RECT 45.785000   0.305000 49.365000   0.375000 ;
      RECT 45.785000   0.375000 49.310000   0.430000 ;
      RECT 45.785000   0.430000 49.310000   1.105000 ;
      RECT 45.785000   1.105000 66.260000   4.865000 ;
      RECT 45.785000   1.105000 66.260000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.240000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   1.755000 67.995000   4.865000 ;
      RECT 45.785000   4.240000 76.870000   4.865000 ;
      RECT 45.855000   4.865000 76.870000   4.935000 ;
      RECT 45.855000   4.865000 76.870000   4.935000 ;
      RECT 45.925000   4.935000 76.870000   5.005000 ;
      RECT 45.925000   4.935000 76.870000   5.005000 ;
      RECT 45.995000   5.005000 76.870000   5.075000 ;
      RECT 45.995000   5.005000 76.870000   5.075000 ;
      RECT 46.065000   5.075000 76.870000   5.145000 ;
      RECT 46.065000   5.075000 76.870000   5.145000 ;
      RECT 46.100000   5.375000 78.570000   5.530000 ;
      RECT 46.135000   5.145000 76.870000   5.215000 ;
      RECT 46.135000   5.145000 76.870000   5.215000 ;
      RECT 46.205000   5.215000 76.870000   5.285000 ;
      RECT 46.205000   5.215000 76.870000   5.285000 ;
      RECT 46.255000   5.530000 78.570000   6.920000 ;
      RECT 46.275000   5.285000 76.870000   5.355000 ;
      RECT 46.275000   5.285000 76.870000   5.355000 ;
      RECT 46.345000   5.355000 76.870000   5.425000 ;
      RECT 46.345000   5.355000 76.870000   5.425000 ;
      RECT 46.395000   5.425000 76.870000   5.475000 ;
      RECT 46.395000   5.425000 76.870000   5.475000 ;
      RECT 46.395000   5.475000 76.870000   5.515000 ;
      RECT 46.395000   5.515000 78.430000   7.060000 ;
      RECT 49.310000   0.000000 49.575000   0.165000 ;
      RECT 50.255000   0.000000 66.695000   0.240000 ;
      RECT 50.255000   0.240000 66.695000   0.485000 ;
      RECT 50.395000   0.000000 50.640000   0.185000 ;
      RECT 50.465000   0.185000 66.555000   0.255000 ;
      RECT 50.500000   0.485000 66.695000   0.840000 ;
      RECT 50.500000   0.840000 66.570000   0.965000 ;
      RECT 50.535000   0.255000 66.555000   0.325000 ;
      RECT 50.605000   0.325000 66.555000   0.395000 ;
      RECT 50.640000   0.000000 66.260000   4.865000 ;
      RECT 50.640000   0.395000 66.555000   0.430000 ;
      RECT 50.640000   0.785000 66.485000   0.855000 ;
      RECT 50.640000   0.855000 66.415000   0.925000 ;
      RECT 50.640000   0.925000 66.345000   0.995000 ;
      RECT 50.640000   0.995000 66.275000   1.065000 ;
      RECT 50.640000   1.065000 66.260000   1.080000 ;
      RECT 66.260000   0.000000 66.555000   0.185000 ;
      RECT 66.260000   0.430000 66.555000   0.785000 ;
      RECT 67.235000   0.000000 68.135000   0.870000 ;
      RECT 67.235000   0.870000 68.135000   1.135000 ;
      RECT 67.375000   0.000000 67.995000   0.815000 ;
      RECT 67.445000   0.815000 67.995000   0.885000 ;
      RECT 67.500000   1.135000 68.135000   1.615000 ;
      RECT 67.515000   0.885000 67.995000   0.955000 ;
      RECT 67.585000   0.955000 67.995000   1.025000 ;
      RECT 67.640000   1.025000 67.995000   1.080000 ;
      RECT 67.640000   1.080000 67.995000   1.755000 ;
      RECT 69.065000   0.000000 76.140000   2.110000 ;
      RECT 69.065000   2.110000 77.010000   2.985000 ;
      RECT 69.065000   2.985000 77.010000   4.100000 ;
      RECT 69.205000   0.000000 76.000000   3.005000 ;
      RECT 69.205000   2.170000 76.000000   2.240000 ;
      RECT 69.205000   2.170000 76.000000   2.240000 ;
      RECT 69.205000   2.240000 76.070000   2.310000 ;
      RECT 69.205000   2.240000 76.070000   2.310000 ;
      RECT 69.205000   2.310000 76.140000   2.380000 ;
      RECT 69.205000   2.310000 76.140000   2.380000 ;
      RECT 69.205000   2.380000 76.210000   2.450000 ;
      RECT 69.205000   2.380000 76.210000   2.450000 ;
      RECT 69.205000   2.450000 76.280000   2.520000 ;
      RECT 69.205000   2.450000 76.280000   2.520000 ;
      RECT 69.205000   2.520000 76.350000   2.590000 ;
      RECT 69.205000   2.520000 76.350000   2.590000 ;
      RECT 69.205000   2.590000 76.420000   2.660000 ;
      RECT 69.205000   2.590000 76.420000   2.660000 ;
      RECT 69.205000   2.660000 76.490000   2.730000 ;
      RECT 69.205000   2.660000 76.490000   2.730000 ;
      RECT 69.205000   2.730000 76.560000   2.800000 ;
      RECT 69.205000   2.730000 76.560000   2.800000 ;
      RECT 69.205000   2.800000 76.630000   2.870000 ;
      RECT 69.205000   2.800000 76.630000   2.870000 ;
      RECT 69.205000   2.870000 76.700000   2.940000 ;
      RECT 69.205000   2.870000 76.700000   2.940000 ;
      RECT 69.205000   2.940000 76.770000   3.010000 ;
      RECT 69.205000   2.940000 76.770000   3.010000 ;
      RECT 69.205000   3.010000 76.840000   3.040000 ;
      RECT 69.205000   3.010000 76.840000   3.040000 ;
      RECT 69.205000   3.040000 76.870000   4.240000 ;
      RECT 76.570000  50.910000 79.435000  52.365000 ;
      RECT 76.570000  52.365000 79.435000  53.050000 ;
      RECT 76.710000  50.965000 79.435000  52.310000 ;
      RECT 76.775000  50.900000 79.435000  50.965000 ;
      RECT 76.780000  52.310000 79.435000  52.380000 ;
      RECT 76.845000  50.830000 79.435000  50.900000 ;
      RECT 76.850000  52.380000 79.435000  52.450000 ;
      RECT 76.915000  50.760000 79.435000  50.830000 ;
      RECT 76.920000  52.450000 79.435000  52.520000 ;
      RECT 76.985000  50.690000 79.435000  50.760000 ;
      RECT 76.990000  52.520000 79.435000  52.590000 ;
      RECT 77.055000  50.620000 79.435000  50.690000 ;
      RECT 77.060000   0.000000 77.470000   0.925000 ;
      RECT 77.060000   0.925000 77.350000   1.045000 ;
      RECT 77.060000   1.045000 77.250000   1.565000 ;
      RECT 77.060000   1.565000 77.250000   1.605000 ;
      RECT 77.060000  52.590000 79.435000  52.660000 ;
      RECT 77.100000   1.605000 78.570000   2.535000 ;
      RECT 77.125000  50.550000 79.435000  50.620000 ;
      RECT 77.130000  52.660000 79.435000  52.730000 ;
      RECT 77.195000  50.480000 79.435000  50.550000 ;
      RECT 77.200000  52.730000 79.435000  52.800000 ;
      RECT 77.255000  53.050000 79.435000  96.135000 ;
      RECT 77.255000  96.135000 79.435000  96.280000 ;
      RECT 77.265000  50.410000 79.435000  50.480000 ;
      RECT 77.270000  52.800000 79.435000  52.870000 ;
      RECT 77.335000  50.340000 79.435000  50.410000 ;
      RECT 77.340000  52.870000 79.435000  52.940000 ;
      RECT 77.395000  52.940000 79.435000  52.995000 ;
      RECT 77.395000  52.995000 79.435000  96.080000 ;
      RECT 77.395000  96.280000 80.000000  96.365000 ;
      RECT 77.405000  50.270000 79.435000  50.340000 ;
      RECT 77.465000  96.080000 79.435000  96.150000 ;
      RECT 77.475000  50.200000 79.435000  50.270000 ;
      RECT 77.505000   1.745000 78.430000   1.815000 ;
      RECT 77.535000  96.150000 79.435000  96.220000 ;
      RECT 77.545000  50.130000 79.435000  50.200000 ;
      RECT 77.575000   1.815000 78.430000   1.885000 ;
      RECT 77.595000  96.220000 79.435000  96.280000 ;
      RECT 77.615000  50.060000 79.435000  50.130000 ;
      RECT 77.645000   1.885000 78.430000   1.955000 ;
      RECT 77.665000  96.280000 80.000000  96.350000 ;
      RECT 77.685000  49.990000 79.435000  50.060000 ;
      RECT 77.715000   1.955000 78.430000   2.025000 ;
      RECT 77.735000  96.350000 80.000000  96.420000 ;
      RECT 77.755000  49.920000 79.435000  49.990000 ;
      RECT 77.785000   2.025000 78.430000   2.095000 ;
      RECT 77.805000  96.420000 80.000000  96.490000 ;
      RECT 77.820000  96.490000 80.000000  96.505000 ;
      RECT 77.825000  49.850000 79.435000  49.920000 ;
      RECT 77.855000   2.095000 78.430000   2.165000 ;
      RECT 77.895000  49.780000 79.435000  49.850000 ;
      RECT 77.925000   2.165000 78.430000   2.235000 ;
      RECT 77.965000  49.710000 79.435000  49.780000 ;
      RECT 77.995000   2.235000 78.430000   2.305000 ;
      RECT 78.010000   0.000000 78.565000   0.815000 ;
      RECT 78.010000   0.815000 78.565000   1.045000 ;
      RECT 78.030000   2.535000 78.570000   5.375000 ;
      RECT 78.035000  49.640000 79.435000  49.710000 ;
      RECT 78.065000   2.305000 78.430000   2.375000 ;
      RECT 78.105000  49.570000 79.435000  49.640000 ;
      RECT 78.135000   2.375000 78.430000   2.445000 ;
      RECT 78.150000   0.000000 78.425000   0.760000 ;
      RECT 78.170000   2.445000 78.430000   2.480000 ;
      RECT 78.170000   2.480000 78.430000   5.515000 ;
      RECT 78.175000  49.500000 79.435000  49.570000 ;
      RECT 78.220000   0.760000 78.425000   0.830000 ;
      RECT 78.245000  49.430000 79.435000  49.500000 ;
      RECT 78.290000   0.830000 78.425000   0.900000 ;
      RECT 78.295000   0.900000 78.425000   0.905000 ;
      RECT 78.315000  49.360000 79.435000  49.430000 ;
      RECT 78.350000   1.045000 78.565000   1.275000 ;
      RECT 78.350000   1.275000 78.570000   1.280000 ;
      RECT 78.350000   1.280000 78.570000   1.605000 ;
      RECT 78.385000  49.290000 79.435000  49.360000 ;
      RECT 78.455000  49.220000 79.435000  49.290000 ;
      RECT 78.525000  49.150000 79.435000  49.220000 ;
      RECT 78.595000  49.080000 79.435000  49.150000 ;
      RECT 78.665000  49.010000 79.435000  49.080000 ;
      RECT 78.735000  48.940000 79.435000  49.010000 ;
      RECT 78.805000  48.870000 79.435000  48.940000 ;
      RECT 78.875000  48.800000 79.435000  48.870000 ;
      RECT 78.945000  10.505000 79.435000  16.185000 ;
      RECT 78.945000  16.185000 79.435000  16.675000 ;
      RECT 78.945000  48.730000 79.435000  48.800000 ;
      RECT 79.015000  48.660000 79.435000  48.730000 ;
      RECT 79.045000   0.000000 79.435000   1.065000 ;
      RECT 79.045000   1.065000 79.435000   1.070000 ;
      RECT 79.050000   1.070000 79.435000  10.400000 ;
      RECT 79.050000  10.400000 79.435000  10.505000 ;
      RECT 79.085000  10.560000 79.435000  16.130000 ;
      RECT 79.085000  48.590000 79.435000  48.660000 ;
      RECT 79.135000  10.510000 79.435000  10.560000 ;
      RECT 79.155000  16.130000 79.435000  16.200000 ;
      RECT 79.155000  48.520000 79.435000  48.590000 ;
      RECT 79.185000   0.000000 79.435000   1.010000 ;
      RECT 79.190000   1.010000 79.435000   1.015000 ;
      RECT 79.190000   1.015000 79.435000  10.455000 ;
      RECT 79.190000  10.455000 79.435000  10.510000 ;
      RECT 79.225000  16.200000 79.435000  16.270000 ;
      RECT 79.225000  48.450000 79.435000  48.520000 ;
      RECT 79.295000  16.270000 79.435000  16.340000 ;
      RECT 79.295000  48.380000 79.435000  48.450000 ;
      RECT 79.365000  16.340000 79.435000  16.410000 ;
      RECT 79.365000  48.310000 79.435000  48.380000 ;
    LAYER met3 ;
      RECT  0.000000   0.000000  0.100000 106.585000 ;
      RECT  0.000000 118.955000  0.100000 178.610000 ;
      RECT  0.000000 178.610000  2.960000 181.470000 ;
      RECT  0.000000 178.800000  0.150000 178.950000 ;
      RECT  0.000000 178.950000  0.300000 179.100000 ;
      RECT  0.000000 179.100000  0.450000 179.250000 ;
      RECT  0.000000 179.250000  0.600000 179.400000 ;
      RECT  0.000000 179.400000  0.750000 179.550000 ;
      RECT  0.000000 179.550000  0.900000 179.700000 ;
      RECT  0.000000 179.700000  1.050000 179.850000 ;
      RECT  0.000000 179.850000  1.200000 180.000000 ;
      RECT  0.000000 180.000000  1.350000 180.150000 ;
      RECT  0.000000 180.150000  1.500000 180.300000 ;
      RECT  0.000000 180.300000  1.650000 180.450000 ;
      RECT  0.000000 180.450000  1.800000 180.600000 ;
      RECT  0.000000 180.600000  1.950000 180.750000 ;
      RECT  0.000000 180.750000  2.100000 180.900000 ;
      RECT  0.000000 180.900000  2.250000 181.050000 ;
      RECT  0.000000 181.050000  2.400000 181.200000 ;
      RECT  0.000000 181.200000  2.550000 181.350000 ;
      RECT  0.000000 181.350000  2.700000 181.500000 ;
      RECT  0.000000 181.470000 80.000000 200.000000 ;
      RECT  0.000000 181.500000  2.850000 181.570000 ;
      RECT  0.000000 181.570000  7.970000 184.570000 ;
      RECT  0.000000 184.570000  7.965000 184.575000 ;
      RECT  0.000000 184.575000  3.005000 196.995000 ;
      RECT  0.000000 196.995000 80.000000 200.000000 ;
      RECT  1.320000   0.000000 45.565000  36.930000 ;
      RECT  1.320000  36.930000 46.275000  37.640000 ;
      RECT  1.320000  37.640000 60.310000  47.660000 ;
      RECT  1.320000  47.660000 61.410000  74.310000 ;
      RECT  1.320000  74.310000 62.735000  75.635000 ;
      RECT  1.320000  75.635000 68.390000  76.345000 ;
      RECT  1.320000  76.345000 68.390000 102.210000 ;
      RECT  1.320000 102.210000 78.280000 106.585000 ;
      RECT  1.320000 118.955000 78.280000 176.780000 ;
      RECT  1.320000 176.780000 80.000000 178.110000 ;
      RECT  1.320000 178.110000 80.000000 180.140000 ;
      RECT  1.415000   0.945000 45.465000   1.675000 ;
      RECT  1.420000   0.000000 45.465000   0.945000 ;
      RECT  1.420000   1.675000 45.465000   3.950000 ;
      RECT  1.420000   3.950000  4.425000  36.970000 ;
      RECT  1.420000  36.970000 45.465000  37.120000 ;
      RECT  1.420000  37.120000 45.615000  37.270000 ;
      RECT  1.420000  37.270000 45.765000  37.420000 ;
      RECT  1.420000  37.420000 45.915000  37.570000 ;
      RECT  1.420000  37.570000 46.065000  37.720000 ;
      RECT  1.420000  37.720000 46.215000  37.740000 ;
      RECT  1.420000  37.740000  4.425000  74.350000 ;
      RECT  1.420000  74.350000 61.310000  74.500000 ;
      RECT  1.420000  74.500000 61.460000  74.650000 ;
      RECT  1.420000  74.650000 61.610000  74.800000 ;
      RECT  1.420000  74.800000 61.760000  74.950000 ;
      RECT  1.420000  74.950000 61.910000  75.100000 ;
      RECT  1.420000  75.100000 62.060000  75.250000 ;
      RECT  1.420000  75.250000 62.210000  75.400000 ;
      RECT  1.420000  75.400000 62.360000  75.550000 ;
      RECT  1.420000  75.550000 62.510000  75.700000 ;
      RECT  1.420000  75.700000 62.660000  75.735000 ;
      RECT  1.420000  75.735000 67.640000  75.885000 ;
      RECT  1.420000  75.885000 67.790000  76.035000 ;
      RECT  1.420000  76.035000 67.940000  76.185000 ;
      RECT  1.420000  76.185000 68.090000  76.335000 ;
      RECT  1.420000  76.335000 68.240000  76.385000 ;
      RECT  1.420000  76.385000 68.290000 106.585000 ;
      RECT  1.420000 118.955000  4.460000 121.960000 ;
      RECT  1.420000 121.960000  4.425000 173.875000 ;
      RECT  1.420000 173.875000  4.475000 176.880000 ;
      RECT  1.420000 176.880000  4.475000 176.960000 ;
      RECT  1.420000 176.960000  4.555000 177.040000 ;
      RECT  1.420000 177.040000  7.970000 178.070000 ;
      RECT  1.440000 178.070000 80.000000 178.090000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 102.310000 78.180000 118.955000 ;
      RECT  1.460000 178.090000 80.000000 178.110000 ;
      RECT  1.460000 178.110000  7.970000 178.145000 ;
      RECT  1.645000 178.145000 80.000000 178.295000 ;
      RECT  1.795000 178.295000 80.000000 178.445000 ;
      RECT  1.945000 178.445000 80.000000 178.595000 ;
      RECT  2.000000 106.585000 78.280000 118.955000 ;
      RECT  2.095000 178.595000 80.000000 178.745000 ;
      RECT  2.245000 178.745000 80.000000 178.895000 ;
      RECT  2.395000 178.895000 80.000000 179.045000 ;
      RECT  2.545000 179.045000 80.000000 179.195000 ;
      RECT  2.695000 179.195000 80.000000 179.345000 ;
      RECT  2.845000 179.345000 80.000000 179.495000 ;
      RECT  2.995000 179.495000 80.000000 179.645000 ;
      RECT  3.000000 184.570000 77.000000 197.000000 ;
      RECT  3.145000 179.645000 80.000000 179.795000 ;
      RECT  3.295000 179.795000 80.000000 179.945000 ;
      RECT  3.390000 179.945000 80.000000 180.040000 ;
      RECT  4.420000   3.000000 42.465000  38.215000 ;
      RECT  4.420000  38.215000 42.465000  38.365000 ;
      RECT  4.420000  38.215000 42.465000  38.365000 ;
      RECT  4.420000  38.365000 42.615000  38.515000 ;
      RECT  4.420000  38.365000 42.615000  38.515000 ;
      RECT  4.420000  38.515000 42.765000  38.665000 ;
      RECT  4.420000  38.515000 42.765000  38.665000 ;
      RECT  4.420000  38.665000 42.915000  38.815000 ;
      RECT  4.420000  38.665000 42.915000  38.815000 ;
      RECT  4.420000  38.815000 43.065000  38.965000 ;
      RECT  4.420000  38.815000 43.065000  38.965000 ;
      RECT  4.420000  38.965000 43.215000  39.115000 ;
      RECT  4.420000  38.965000 43.215000  39.115000 ;
      RECT  4.420000  39.115000 43.365000  39.265000 ;
      RECT  4.420000  39.115000 43.365000  39.265000 ;
      RECT  4.420000  39.265000 43.515000  39.415000 ;
      RECT  4.420000  39.265000 43.515000  39.415000 ;
      RECT  4.420000  39.415000 43.665000  39.565000 ;
      RECT  4.420000  39.415000 43.665000  39.565000 ;
      RECT  4.420000  39.565000 43.815000  39.715000 ;
      RECT  4.420000  39.565000 43.815000  39.715000 ;
      RECT  4.420000  39.715000 43.965000  39.865000 ;
      RECT  4.420000  39.715000 43.965000  39.865000 ;
      RECT  4.420000  39.865000 44.115000  40.015000 ;
      RECT  4.420000  39.865000 44.115000  40.015000 ;
      RECT  4.420000  40.015000 44.265000  40.165000 ;
      RECT  4.420000  40.015000 44.265000  40.165000 ;
      RECT  4.420000  40.165000 44.415000  40.315000 ;
      RECT  4.420000  40.165000 44.415000  40.315000 ;
      RECT  4.420000  40.315000 44.565000  40.465000 ;
      RECT  4.420000  40.315000 44.565000  40.465000 ;
      RECT  4.420000  40.465000 44.715000  40.615000 ;
      RECT  4.420000  40.465000 44.715000  40.615000 ;
      RECT  4.420000  40.615000 44.865000  40.740000 ;
      RECT  4.420000  40.615000 44.865000  40.740000 ;
      RECT  4.420000  40.740000 57.210000  50.760000 ;
      RECT  4.420000  50.760000 58.310000  75.595000 ;
      RECT  4.420000  75.595000 58.310000  75.745000 ;
      RECT  4.420000  75.595000 58.310000  75.745000 ;
      RECT  4.420000  75.745000 58.460000  75.895000 ;
      RECT  4.420000  75.745000 58.460000  75.895000 ;
      RECT  4.420000  75.895000 58.610000  76.045000 ;
      RECT  4.420000  75.895000 58.610000  76.045000 ;
      RECT  4.420000  76.045000 58.760000  76.195000 ;
      RECT  4.420000  76.045000 58.760000  76.195000 ;
      RECT  4.420000  76.195000 58.910000  76.345000 ;
      RECT  4.420000  76.195000 58.910000  76.345000 ;
      RECT  4.420000  76.345000 59.060000  76.495000 ;
      RECT  4.420000  76.345000 59.060000  76.495000 ;
      RECT  4.420000  76.495000 59.210000  76.645000 ;
      RECT  4.420000  76.495000 59.210000  76.645000 ;
      RECT  4.420000  76.645000 59.360000  76.795000 ;
      RECT  4.420000  76.645000 59.360000  76.795000 ;
      RECT  4.420000  76.795000 59.510000  76.945000 ;
      RECT  4.420000  76.795000 59.510000  76.945000 ;
      RECT  4.420000  76.945000 59.660000  77.095000 ;
      RECT  4.420000  76.945000 59.660000  77.095000 ;
      RECT  4.420000  77.095000 59.810000  77.245000 ;
      RECT  4.420000  77.095000 59.810000  77.245000 ;
      RECT  4.420000  77.245000 59.960000  77.395000 ;
      RECT  4.420000  77.245000 59.960000  77.395000 ;
      RECT  4.420000  77.395000 60.110000  77.545000 ;
      RECT  4.420000  77.395000 60.110000  77.545000 ;
      RECT  4.420000  77.545000 60.260000  77.695000 ;
      RECT  4.420000  77.545000 60.260000  77.695000 ;
      RECT  4.420000  77.695000 60.410000  77.845000 ;
      RECT  4.420000  77.695000 60.410000  77.845000 ;
      RECT  4.420000  77.845000 60.560000  77.995000 ;
      RECT  4.420000  77.845000 60.560000  77.995000 ;
      RECT  4.420000  77.995000 60.710000  78.145000 ;
      RECT  4.420000  77.995000 60.710000  78.145000 ;
      RECT  4.420000  78.145000 60.860000  78.295000 ;
      RECT  4.420000  78.145000 60.860000  78.295000 ;
      RECT  4.420000  78.295000 61.010000  78.445000 ;
      RECT  4.420000  78.295000 61.010000  78.445000 ;
      RECT  4.420000  78.445000 61.160000  78.595000 ;
      RECT  4.420000  78.445000 61.160000  78.595000 ;
      RECT  4.420000  78.595000 61.310000  78.735000 ;
      RECT  4.420000  78.595000 61.310000  78.735000 ;
      RECT  4.420000  78.735000 65.285000 103.585000 ;
      RECT  4.420000 121.955000 75.175000 176.825000 ;
      RECT  4.460000 103.585000 65.285000 105.310000 ;
      RECT  4.460000 105.310000 75.175000 121.955000 ;
      RECT  4.525000 176.825000 75.175000 176.930000 ;
      RECT  4.525000 176.825000 75.175000 176.930000 ;
      RECT  4.630000 176.930000 75.175000 177.035000 ;
      RECT  4.630000 176.930000 75.175000 177.035000 ;
      RECT  4.635000 177.035000 75.175000 177.040000 ;
      RECT  4.635000 177.035000 75.175000 177.040000 ;
      RECT  4.865000 180.140000 80.000000 181.470000 ;
      RECT  4.965000 178.070000  7.970000 178.110000 ;
      RECT  4.965000 178.145000  7.970000 181.570000 ;
      RECT  7.965000 177.040000 75.175000 179.880000 ;
      RECT  7.965000 179.880000 77.000000 184.570000 ;
      RECT 42.460000   3.950000 45.465000  36.970000 ;
      RECT 42.465000  37.740000 52.000000  40.745000 ;
      RECT 46.495000   0.000000 62.520000   5.430000 ;
      RECT 46.495000   5.430000 61.960000   5.990000 ;
      RECT 46.495000   5.990000 59.300000   7.300000 ;
      RECT 46.495000   7.300000 59.300000  11.060000 ;
      RECT 46.495000  11.060000 61.170000  12.930000 ;
      RECT 46.495000  12.930000 61.170000  18.080000 ;
      RECT 46.495000  18.080000 60.310000  18.940000 ;
      RECT 46.495000  18.940000 60.310000  35.570000 ;
      RECT 46.495000  35.570000 47.660000  36.315000 ;
      RECT 46.495000  36.315000 47.880000  36.535000 ;
      RECT 46.495000  36.535000 47.880000  36.540000 ;
      RECT 46.495000  36.540000 47.880000  36.610000 ;
      RECT 46.565000  36.610000 47.780000  36.710000 ;
      RECT 46.595000   0.000000 62.420000   3.005000 ;
      RECT 46.595000   3.005000 49.600000   5.390000 ;
      RECT 46.595000   5.390000 62.270000   5.540000 ;
      RECT 46.595000   5.540000 62.120000   5.690000 ;
      RECT 46.595000   5.690000 61.970000   5.840000 ;
      RECT 46.595000   5.840000 61.920000   5.890000 ;
      RECT 46.595000   5.890000 60.420000   6.040000 ;
      RECT 46.595000   6.040000 60.270000   6.190000 ;
      RECT 46.595000   6.190000 60.120000   6.340000 ;
      RECT 46.595000   6.340000 59.970000   6.490000 ;
      RECT 46.595000   6.490000 59.820000   6.640000 ;
      RECT 46.595000   6.640000 59.670000   6.790000 ;
      RECT 46.595000   6.790000 59.520000   6.940000 ;
      RECT 46.595000   6.940000 59.370000   7.090000 ;
      RECT 46.595000   7.090000 59.220000   7.240000 ;
      RECT 46.595000   7.240000 59.200000   7.260000 ;
      RECT 46.595000   7.260000 59.200000  35.470000 ;
      RECT 46.595000  11.100000 59.200000  11.250000 ;
      RECT 46.595000  11.250000 59.350000  11.400000 ;
      RECT 46.595000  11.400000 59.500000  11.550000 ;
      RECT 46.595000  11.550000 59.650000  11.700000 ;
      RECT 46.595000  11.700000 59.800000  11.850000 ;
      RECT 46.595000  11.850000 59.950000  12.000000 ;
      RECT 46.595000  12.000000 60.100000  12.150000 ;
      RECT 46.595000  12.150000 60.250000  12.300000 ;
      RECT 46.595000  12.300000 60.400000  12.450000 ;
      RECT 46.595000  12.450000 60.550000  12.600000 ;
      RECT 46.595000  12.600000 60.700000  12.750000 ;
      RECT 46.595000  12.750000 60.850000  12.900000 ;
      RECT 46.595000  12.900000 61.000000  12.970000 ;
      RECT 46.595000  18.040000 60.920000  18.190000 ;
      RECT 46.595000  18.190000 60.770000  18.340000 ;
      RECT 46.595000  18.340000 60.620000  18.490000 ;
      RECT 46.595000  18.490000 60.470000  18.640000 ;
      RECT 46.595000  18.640000 60.320000  18.790000 ;
      RECT 46.595000  18.790000 60.210000  18.900000 ;
      RECT 46.595000  35.470000 47.560000  36.355000 ;
      RECT 46.595000  36.355000 47.560000  36.425000 ;
      RECT 46.595000  36.425000 47.630000  36.495000 ;
      RECT 46.595000  36.495000 47.700000  36.500000 ;
      RECT 46.650000  36.500000 47.705000  36.555000 ;
      RECT 46.705000  36.555000 47.760000  36.610000 ;
      RECT 48.310000  37.640000 60.210000  37.740000 ;
      RECT 48.460000  37.490000 60.210000  37.640000 ;
      RECT 48.610000  37.340000 60.210000  37.490000 ;
      RECT 48.760000  37.190000 60.210000  37.340000 ;
      RECT 48.810000  36.545000 60.310000  37.000000 ;
      RECT 48.810000  37.000000 60.310000  37.640000 ;
      RECT 48.910000  36.585000 52.145000  37.040000 ;
      RECT 48.910000  37.040000 60.210000  37.190000 ;
      RECT 49.025000  36.470000 60.210000  36.585000 ;
      RECT 49.040000  35.570000 60.310000  36.315000 ;
      RECT 49.040000  36.315000 60.310000  36.545000 ;
      RECT 49.140000  35.470000 52.145000  36.585000 ;
      RECT 49.140000  36.355000 60.210000  36.470000 ;
      RECT 49.510000  40.685000 57.210000  40.740000 ;
      RECT 49.510000  40.685000 57.210000  40.740000 ;
      RECT 49.595000   3.000000 59.065000   3.150000 ;
      RECT 49.595000   3.000000 59.065000   3.150000 ;
      RECT 49.595000   3.150000 58.915000   3.300000 ;
      RECT 49.595000   3.150000 58.915000   3.300000 ;
      RECT 49.595000   3.300000 58.765000   3.450000 ;
      RECT 49.595000   3.300000 58.765000   3.450000 ;
      RECT 49.595000   3.450000 58.615000   3.600000 ;
      RECT 49.595000   3.450000 58.615000   3.600000 ;
      RECT 49.595000   3.600000 58.465000   3.750000 ;
      RECT 49.595000   3.600000 58.465000   3.750000 ;
      RECT 49.595000   3.750000 58.315000   3.900000 ;
      RECT 49.595000   3.750000 58.315000   3.900000 ;
      RECT 49.595000   3.900000 58.165000   4.050000 ;
      RECT 49.595000   3.900000 58.165000   4.050000 ;
      RECT 49.595000   4.050000 58.015000   4.200000 ;
      RECT 49.595000   4.050000 58.015000   4.200000 ;
      RECT 49.595000   4.200000 57.865000   4.350000 ;
      RECT 49.595000   4.200000 57.865000   4.350000 ;
      RECT 49.595000   4.350000 57.715000   4.500000 ;
      RECT 49.595000   4.350000 57.715000   4.500000 ;
      RECT 49.595000   4.500000 57.565000   4.650000 ;
      RECT 49.595000   4.500000 57.565000   4.650000 ;
      RECT 49.595000   4.650000 57.415000   4.800000 ;
      RECT 49.595000   4.650000 57.415000   4.800000 ;
      RECT 49.595000   4.800000 57.265000   4.950000 ;
      RECT 49.595000   4.800000 57.265000   4.950000 ;
      RECT 49.595000   4.950000 57.115000   5.100000 ;
      RECT 49.595000   4.950000 57.115000   5.100000 ;
      RECT 49.595000   5.100000 56.965000   5.250000 ;
      RECT 49.595000   5.100000 56.965000   5.250000 ;
      RECT 49.595000   5.250000 56.815000   5.400000 ;
      RECT 49.595000   5.250000 56.815000   5.400000 ;
      RECT 49.595000   5.400000 56.665000   5.550000 ;
      RECT 49.595000   5.400000 56.665000   5.550000 ;
      RECT 49.595000   5.550000 56.515000   5.700000 ;
      RECT 49.595000   5.550000 56.515000   5.700000 ;
      RECT 49.595000   5.700000 56.365000   5.850000 ;
      RECT 49.595000   5.700000 56.365000   5.850000 ;
      RECT 49.595000   5.850000 56.215000   6.000000 ;
      RECT 49.595000   5.850000 56.215000   6.000000 ;
      RECT 49.595000   6.000000 56.200000   6.015000 ;
      RECT 49.595000   6.000000 56.200000   6.015000 ;
      RECT 49.595000   6.015000 56.200000  12.345000 ;
      RECT 49.595000  12.345000 56.200000  12.495000 ;
      RECT 49.595000  12.345000 56.200000  12.495000 ;
      RECT 49.595000  12.495000 56.350000  12.645000 ;
      RECT 49.595000  12.495000 56.350000  12.645000 ;
      RECT 49.595000  12.645000 56.500000  12.795000 ;
      RECT 49.595000  12.645000 56.500000  12.795000 ;
      RECT 49.595000  12.795000 56.650000  12.945000 ;
      RECT 49.595000  12.795000 56.650000  12.945000 ;
      RECT 49.595000  12.945000 56.800000  13.095000 ;
      RECT 49.595000  12.945000 56.800000  13.095000 ;
      RECT 49.595000  13.095000 56.950000  13.245000 ;
      RECT 49.595000  13.095000 56.950000  13.245000 ;
      RECT 49.595000  13.245000 57.100000  13.395000 ;
      RECT 49.595000  13.245000 57.100000  13.395000 ;
      RECT 49.595000  13.395000 57.250000  13.545000 ;
      RECT 49.595000  13.395000 57.250000  13.545000 ;
      RECT 49.595000  13.545000 57.400000  13.695000 ;
      RECT 49.595000  13.545000 57.400000  13.695000 ;
      RECT 49.595000  13.695000 57.550000  13.845000 ;
      RECT 49.595000  13.695000 57.550000  13.845000 ;
      RECT 49.595000  13.845000 57.700000  13.995000 ;
      RECT 49.595000  13.845000 57.700000  13.995000 ;
      RECT 49.595000  13.995000 57.850000  14.145000 ;
      RECT 49.595000  13.995000 57.850000  14.145000 ;
      RECT 49.595000  14.145000 58.000000  14.215000 ;
      RECT 49.595000  14.145000 58.000000  14.215000 ;
      RECT 49.595000  14.215000 58.070000  16.795000 ;
      RECT 49.595000  16.795000 57.920000  16.945000 ;
      RECT 49.595000  16.795000 57.920000  16.945000 ;
      RECT 49.595000  16.945000 57.770000  17.095000 ;
      RECT 49.595000  16.945000 57.770000  17.095000 ;
      RECT 49.595000  17.095000 57.620000  17.245000 ;
      RECT 49.595000  17.095000 57.620000  17.245000 ;
      RECT 49.595000  17.245000 57.470000  17.395000 ;
      RECT 49.595000  17.245000 57.470000  17.395000 ;
      RECT 49.595000  17.395000 57.320000  17.545000 ;
      RECT 49.595000  17.395000 57.320000  17.545000 ;
      RECT 49.595000  17.545000 57.210000  17.655000 ;
      RECT 49.595000  17.545000 57.210000  17.655000 ;
      RECT 49.595000  17.655000 57.210000  32.470000 ;
      RECT 49.660000  40.535000 57.210000  40.685000 ;
      RECT 49.660000  40.535000 57.210000  40.685000 ;
      RECT 49.810000  40.385000 57.210000  40.535000 ;
      RECT 49.810000  40.385000 57.210000  40.535000 ;
      RECT 49.960000  40.235000 57.210000  40.385000 ;
      RECT 49.960000  40.235000 57.210000  40.385000 ;
      RECT 50.110000  40.085000 57.210000  40.235000 ;
      RECT 50.110000  40.085000 57.210000  40.235000 ;
      RECT 50.260000  39.935000 57.210000  40.085000 ;
      RECT 50.260000  39.935000 57.210000  40.085000 ;
      RECT 50.410000  39.785000 57.210000  39.935000 ;
      RECT 50.410000  39.785000 57.210000  39.935000 ;
      RECT 50.560000  39.635000 57.210000  39.785000 ;
      RECT 50.560000  39.635000 57.210000  39.785000 ;
      RECT 50.710000  39.485000 57.210000  39.635000 ;
      RECT 50.710000  39.485000 57.210000  39.635000 ;
      RECT 50.860000  39.335000 57.210000  39.485000 ;
      RECT 50.860000  39.335000 57.210000  39.485000 ;
      RECT 51.010000  39.185000 57.210000  39.335000 ;
      RECT 51.010000  39.185000 57.210000  39.335000 ;
      RECT 51.160000  39.035000 57.210000  39.185000 ;
      RECT 51.160000  39.035000 57.210000  39.185000 ;
      RECT 51.310000  38.885000 57.210000  39.035000 ;
      RECT 51.310000  38.885000 57.210000  39.035000 ;
      RECT 51.460000  38.735000 57.210000  38.885000 ;
      RECT 51.460000  38.735000 57.210000  38.885000 ;
      RECT 51.610000  38.585000 57.210000  38.735000 ;
      RECT 51.610000  38.585000 57.210000  38.735000 ;
      RECT 51.760000  38.435000 57.210000  38.585000 ;
      RECT 51.760000  38.435000 57.210000  38.585000 ;
      RECT 51.910000  37.830000 57.210000  38.285000 ;
      RECT 51.910000  38.285000 57.210000  38.435000 ;
      RECT 51.910000  38.285000 57.210000  38.435000 ;
      RECT 52.025000  37.715000 57.210000  37.830000 ;
      RECT 52.025000  37.715000 57.210000  37.830000 ;
      RECT 52.140000  32.470000 57.210000  37.600000 ;
      RECT 52.140000  37.600000 57.210000  37.715000 ;
      RECT 52.140000  37.600000 57.210000  37.715000 ;
      RECT 56.825000   3.005000 62.420000   5.390000 ;
      RECT 57.205000  18.900000 60.210000  37.040000 ;
      RECT 57.205000  37.740000 60.210000  47.760000 ;
      RECT 57.210000  47.760000 61.310000  50.765000 ;
      RECT 58.065000  12.970000 61.070000  18.040000 ;
      RECT 58.305000  50.765000 61.310000  74.350000 ;
      RECT 60.685000   7.875000 62.520000   7.930000 ;
      RECT 60.685000   7.930000 62.520000  10.485000 ;
      RECT 60.685000  10.485000 62.520000  12.320000 ;
      RECT 60.785000   7.915000 62.365000   7.945000 ;
      RECT 60.785000   7.945000 62.395000   7.970000 ;
      RECT 60.785000   7.970000 62.420000  10.445000 ;
      RECT 60.930000   7.770000 62.220000   7.915000 ;
      RECT 60.935000  10.445000 62.420000  10.595000 ;
      RECT 61.080000   7.620000 62.070000   7.770000 ;
      RECT 61.085000  10.595000 62.420000  10.745000 ;
      RECT 61.190000   7.370000 62.465000   7.875000 ;
      RECT 61.230000   7.470000 61.920000   7.620000 ;
      RECT 61.235000  10.745000 62.420000  10.895000 ;
      RECT 61.385000  10.895000 62.420000  11.045000 ;
      RECT 61.535000  11.045000 62.420000  11.195000 ;
      RECT 61.685000  11.195000 62.420000  11.345000 ;
      RECT 61.695000  19.515000 62.325000  34.720000 ;
      RECT 61.795000  19.555000 62.225000  34.680000 ;
      RECT 61.795000  34.680000 62.075000  34.830000 ;
      RECT 61.795000  34.830000 61.925000  34.980000 ;
      RECT 61.835000  11.345000 62.420000  11.495000 ;
      RECT 61.925000  19.425000 62.225000  19.555000 ;
      RECT 61.985000  11.495000 62.420000  11.645000 ;
      RECT 62.075000  19.275000 62.225000  19.425000 ;
      RECT 62.135000  11.645000 62.420000  11.795000 ;
      RECT 62.285000  11.795000 62.420000  11.945000 ;
      RECT 63.080000  36.325000 78.280000  72.880000 ;
      RECT 63.080000  72.880000 78.280000  73.965000 ;
      RECT 63.180000  36.365000 67.095000  39.370000 ;
      RECT 63.180000  39.370000 66.185000  69.835000 ;
      RECT 63.180000  69.835000 71.940000  72.840000 ;
      RECT 63.195000  36.350000 78.180000  36.365000 ;
      RECT 63.330000  72.840000 78.180000  72.990000 ;
      RECT 63.345000  36.200000 78.180000  36.350000 ;
      RECT 63.480000  72.990000 78.180000  73.140000 ;
      RECT 63.495000  36.050000 78.180000  36.200000 ;
      RECT 63.630000  73.140000 78.180000  73.290000 ;
      RECT 63.645000  35.900000 78.180000  36.050000 ;
      RECT 63.780000  73.290000 78.180000  73.440000 ;
      RECT 63.795000  35.750000 78.180000  35.900000 ;
      RECT 63.930000  73.440000 78.180000  73.590000 ;
      RECT 63.945000  35.600000 78.180000  35.750000 ;
      RECT 63.995000  18.390000 78.280000  35.410000 ;
      RECT 63.995000  35.410000 78.280000  36.325000 ;
      RECT 64.080000  73.590000 78.180000  73.740000 ;
      RECT 64.095000  18.430000 67.290000  21.435000 ;
      RECT 64.095000  21.435000 67.100000  35.450000 ;
      RECT 64.095000  35.450000 78.180000  35.600000 ;
      RECT 64.190000   0.000000 78.280000  18.195000 ;
      RECT 64.190000  18.195000 78.280000  18.390000 ;
      RECT 64.190000  18.335000 78.180000  18.430000 ;
      RECT 64.205000  73.740000 78.180000  73.865000 ;
      RECT 64.290000   0.000000 78.180000   7.455000 ;
      RECT 64.290000   2.690000 78.180000   2.735000 ;
      RECT 64.290000   2.735000 78.225000   2.780000 ;
      RECT 64.290000   2.780000 78.270000   2.785000 ;
      RECT 64.290000   2.785000 78.180000  18.235000 ;
      RECT 64.290000  18.235000 78.180000  18.335000 ;
      RECT 66.180000  37.610000 75.175000  70.865000 ;
      RECT 66.195000  37.595000 75.175000  37.610000 ;
      RECT 66.195000  37.595000 75.175000  37.610000 ;
      RECT 66.345000  37.445000 75.175000  37.595000 ;
      RECT 66.345000  37.445000 75.175000  37.595000 ;
      RECT 66.495000  37.295000 75.175000  37.445000 ;
      RECT 66.495000  37.295000 75.175000  37.445000 ;
      RECT 66.645000  37.145000 75.175000  37.295000 ;
      RECT 66.645000  37.145000 75.175000  37.295000 ;
      RECT 66.795000  36.995000 75.175000  37.145000 ;
      RECT 66.795000  36.995000 75.175000  37.145000 ;
      RECT 66.945000  36.845000 75.175000  36.995000 ;
      RECT 66.945000  36.845000 75.175000  36.995000 ;
      RECT 67.095000  19.675000 75.175000  36.695000 ;
      RECT 67.095000  36.695000 75.175000  36.845000 ;
      RECT 67.095000  36.695000 75.175000  36.845000 ;
      RECT 67.100000  19.670000 75.175000  19.675000 ;
      RECT 67.100000  19.670000 75.175000  19.675000 ;
      RECT 67.195000  19.575000 75.175000  19.670000 ;
      RECT 67.195000  19.575000 75.175000  19.670000 ;
      RECT 67.290000   3.000000 75.175000   3.935000 ;
      RECT 67.290000   3.935000 75.175000   3.980000 ;
      RECT 67.290000   3.935000 75.175000   3.980000 ;
      RECT 67.290000   3.980000 75.225000   4.025000 ;
      RECT 67.290000   3.980000 75.225000   4.025000 ;
      RECT 67.290000   4.025000 75.270000   4.030000 ;
      RECT 67.290000   4.025000 75.270000   4.030000 ;
      RECT 67.290000   4.030000 75.270000   4.455000 ;
      RECT 67.290000   4.455000 75.175000  19.480000 ;
      RECT 67.290000  19.480000 75.175000  19.575000 ;
      RECT 67.290000  19.480000 75.175000  19.575000 ;
      RECT 68.680000  73.965000 78.280000  75.345000 ;
      RECT 68.870000  73.865000 78.180000  74.015000 ;
      RECT 69.020000  74.015000 78.180000  74.165000 ;
      RECT 69.170000  74.165000 78.180000  74.315000 ;
      RECT 69.320000  74.315000 78.180000  74.465000 ;
      RECT 69.470000  74.465000 78.180000  74.615000 ;
      RECT 69.620000  74.615000 78.180000  74.765000 ;
      RECT 69.770000  74.765000 78.180000  74.915000 ;
      RECT 69.920000  74.915000 78.180000  75.065000 ;
      RECT 70.060000  75.345000 78.280000 102.210000 ;
      RECT 70.070000  75.065000 78.180000  75.215000 ;
      RECT 70.110000  70.865000 75.175000  71.010000 ;
      RECT 70.110000  70.865000 75.175000  71.010000 ;
      RECT 70.160000  73.865000 78.180000 118.955000 ;
      RECT 70.160000  75.215000 78.180000  75.305000 ;
      RECT 70.260000  71.010000 75.175000  71.160000 ;
      RECT 70.260000  71.010000 75.175000  71.160000 ;
      RECT 70.410000  71.160000 75.175000  71.310000 ;
      RECT 70.410000  71.160000 75.175000  71.310000 ;
      RECT 70.560000  71.310000 75.175000  71.460000 ;
      RECT 70.560000  71.310000 75.175000  71.460000 ;
      RECT 70.710000  71.460000 75.175000  71.610000 ;
      RECT 70.710000  71.460000 75.175000  71.610000 ;
      RECT 70.860000  71.610000 75.175000  71.760000 ;
      RECT 70.860000  71.610000 75.175000  71.760000 ;
      RECT 71.010000  71.760000 75.175000  71.910000 ;
      RECT 71.010000  71.760000 75.175000  71.910000 ;
      RECT 71.160000  71.910000 75.175000  72.060000 ;
      RECT 71.160000  71.910000 75.175000  72.060000 ;
      RECT 71.310000  72.060000 75.175000  72.210000 ;
      RECT 71.310000  72.060000 75.175000  72.210000 ;
      RECT 71.460000  72.210000 75.175000  72.360000 ;
      RECT 71.460000  72.210000 75.175000  72.360000 ;
      RECT 71.610000  72.360000 75.175000  72.510000 ;
      RECT 71.610000  72.360000 75.175000  72.510000 ;
      RECT 71.760000  72.510000 75.175000  72.660000 ;
      RECT 71.760000  72.510000 75.175000  72.660000 ;
      RECT 71.910000  72.660000 75.175000  72.810000 ;
      RECT 71.910000  72.660000 75.175000  72.810000 ;
      RECT 72.060000  72.810000 75.175000  72.960000 ;
      RECT 72.060000  72.810000 75.175000  72.960000 ;
      RECT 72.210000  72.960000 75.175000  73.110000 ;
      RECT 72.210000  72.960000 75.175000  73.110000 ;
      RECT 72.360000  73.110000 75.175000  73.260000 ;
      RECT 72.360000  73.110000 75.175000  73.260000 ;
      RECT 72.510000  73.260000 75.175000  73.410000 ;
      RECT 72.510000  73.260000 75.175000  73.410000 ;
      RECT 72.660000  73.410000 75.175000  73.560000 ;
      RECT 72.660000  73.410000 75.175000  73.560000 ;
      RECT 72.810000  73.560000 75.175000  73.710000 ;
      RECT 72.810000  73.560000 75.175000  73.710000 ;
      RECT 72.960000  73.710000 75.175000  73.860000 ;
      RECT 72.960000  73.710000 75.175000  73.860000 ;
      RECT 73.110000  73.860000 75.175000  74.010000 ;
      RECT 73.110000  73.860000 75.175000  74.010000 ;
      RECT 73.160000  74.010000 75.175000  74.060000 ;
      RECT 73.160000  74.010000 75.175000  74.060000 ;
      RECT 73.160000  74.060000 75.175000 105.310000 ;
      RECT 75.175000  18.430000 78.180000  35.450000 ;
      RECT 75.175000  36.365000 78.180000  72.840000 ;
      RECT 75.175000 118.955000 78.180000 176.880000 ;
      RECT 75.175000 176.880000 80.000000 179.885000 ;
      RECT 75.270000   2.785000 78.275000   7.455000 ;
      RECT 76.995000 179.885000 80.000000 196.995000 ;
      RECT 78.180000   1.160000 78.190000   1.490000 ;
      RECT 79.870000   0.000000 80.000000 176.780000 ;
    LAYER met4 ;
      RECT  0.000000   0.000000 80.000000   1.635000 ;
      RECT  0.000000   7.885000  4.675000   8.485000 ;
      RECT  0.000000   7.885000 80.000000   8.485000 ;
      RECT  0.000000  13.935000  4.675000  14.535000 ;
      RECT  0.000000  13.935000 80.000000  14.535000 ;
      RECT  0.000000  18.785000  4.675000  19.385000 ;
      RECT  0.000000  18.785000 80.000000  19.385000 ;
      RECT  0.000000  24.835000  4.675000  25.435000 ;
      RECT  0.000000  24.835000 80.000000  25.435000 ;
      RECT  0.000000  30.885000  4.675000  31.485000 ;
      RECT  0.000000  30.885000 80.000000  31.485000 ;
      RECT  0.000000  35.735000  4.675000  36.335000 ;
      RECT  0.000000  35.735000 80.000000  36.335000 ;
      RECT  0.000000  40.585000  4.675000  41.185000 ;
      RECT  0.000000  40.585000 80.000000  41.185000 ;
      RECT  0.000000  46.635000  4.675000  47.335000 ;
      RECT  0.000000  46.635000 80.000000  47.435000 ;
      RECT  0.000000  57.035000 80.000000  57.835000 ;
      RECT  0.000000  57.135000  4.675000  57.835000 ;
      RECT  0.000000  63.085000  4.675000  63.685000 ;
      RECT  0.000000  63.085000 80.000000  63.685000 ;
      RECT  0.000000  68.935000  4.675000  69.635000 ;
      RECT  0.000000  68.935000 80.000000  69.635000 ;
      RECT  0.000000  95.400000  3.005000 104.215000 ;
      RECT  0.000000  95.400000 80.000000 104.315000 ;
      RECT  0.000000 104.215000  9.485000 104.365000 ;
      RECT  0.000000 104.315000  7.705000 106.285000 ;
      RECT  0.000000 104.365000  9.335000 104.515000 ;
      RECT  0.000000 104.515000  9.185000 104.665000 ;
      RECT  0.000000 104.665000  9.035000 104.815000 ;
      RECT  0.000000 104.815000  8.885000 104.965000 ;
      RECT  0.000000 104.965000  8.735000 105.115000 ;
      RECT  0.000000 105.115000  8.585000 105.265000 ;
      RECT  0.000000 105.265000  8.435000 105.415000 ;
      RECT  0.000000 105.415000  8.285000 105.565000 ;
      RECT  0.000000 105.565000  8.135000 105.715000 ;
      RECT  0.000000 105.715000  7.985000 105.865000 ;
      RECT  0.000000 105.865000  7.835000 106.015000 ;
      RECT  0.000000 106.015000  7.685000 106.165000 ;
      RECT  0.000000 106.165000  7.665000 106.185000 ;
      RECT  0.000000 106.185000  1.600000 106.585000 ;
      RECT  0.000000 106.285000  1.700000 106.585000 ;
      RECT  0.000000 118.955000  1.600000 119.355000 ;
      RECT  0.000000 118.955000  1.700000 119.255000 ;
      RECT  0.000000 119.255000  9.685000 121.550000 ;
      RECT  0.000000 119.355000  7.350000 119.505000 ;
      RECT  0.000000 119.505000  7.500000 119.655000 ;
      RECT  0.000000 119.655000  7.650000 119.805000 ;
      RECT  0.000000 119.805000  7.800000 119.955000 ;
      RECT  0.000000 119.955000  7.950000 120.105000 ;
      RECT  0.000000 120.105000  8.100000 120.255000 ;
      RECT  0.000000 120.255000  8.250000 120.405000 ;
      RECT  0.000000 120.405000  8.400000 120.555000 ;
      RECT  0.000000 120.555000  8.550000 120.705000 ;
      RECT  0.000000 120.705000  8.700000 120.855000 ;
      RECT  0.000000 120.855000  8.850000 121.005000 ;
      RECT  0.000000 121.005000  9.000000 121.155000 ;
      RECT  0.000000 121.155000  9.150000 121.305000 ;
      RECT  0.000000 121.305000  9.300000 121.455000 ;
      RECT  0.000000 121.455000  9.450000 121.605000 ;
      RECT  0.000000 121.550000 80.000000 175.385000 ;
      RECT  0.000000 121.605000  9.600000 121.650000 ;
      RECT  0.000000 121.650000 15.900000 124.655000 ;
      RECT  0.000000 124.655000  3.005000 172.380000 ;
      RECT  0.000000 172.380000  4.670000 175.385000 ;
      RECT  1.365000  14.535000  4.675000  18.785000 ;
      RECT  1.365000  14.535000 78.635000  18.785000 ;
      RECT  1.455000  70.310000  4.675000  94.885000 ;
      RECT  1.570000  47.435000 78.430000  57.035000 ;
      RECT  1.670000   1.635000 78.330000   4.640000 ;
      RECT  1.670000   1.635000 78.330000   7.885000 ;
      RECT  1.670000   4.640000  4.675000   7.885000 ;
      RECT  1.670000   8.485000  4.675000  13.935000 ;
      RECT  1.670000   8.485000 78.330000  13.935000 ;
      RECT  1.670000  19.385000  4.675000  24.835000 ;
      RECT  1.670000  19.385000 78.330000  24.835000 ;
      RECT  1.670000  25.435000  4.675000  30.885000 ;
      RECT  1.670000  25.435000 78.330000  30.885000 ;
      RECT  1.670000  31.485000  4.675000  35.735000 ;
      RECT  1.670000  31.485000 78.330000  35.735000 ;
      RECT  1.670000  36.335000  4.675000  40.585000 ;
      RECT  1.670000  36.335000 78.330000  40.585000 ;
      RECT  1.670000  41.185000  4.675000  46.635000 ;
      RECT  1.670000  41.185000 78.330000  46.635000 ;
      RECT  1.670000  47.335000  4.675000  57.135000 ;
      RECT  1.670000  57.835000  4.675000  63.085000 ;
      RECT  1.670000  57.835000 78.330000  63.085000 ;
      RECT  1.670000  63.685000  4.675000  68.935000 ;
      RECT  1.670000  63.685000 78.330000  68.935000 ;
      RECT  1.670000  69.635000  4.675000  70.310000 ;
      RECT  1.670000  69.635000 78.330000  95.400000 ;
      RECT  1.670000  94.885000 78.330000 104.215000 ;
      RECT  1.670000 175.385000  4.675000 196.995000 ;
      RECT  1.670000 175.385000 78.330000 200.000000 ;
      RECT  1.670000 196.995000 78.330000 200.000000 ;
      RECT  3.000000  98.400000 77.000000 101.210000 ;
      RECT  3.000000 101.210000  8.245000 101.360000 ;
      RECT  3.000000 101.210000  8.245000 101.360000 ;
      RECT  3.000000 101.360000  8.095000 101.510000 ;
      RECT  3.000000 101.360000  8.095000 101.510000 ;
      RECT  3.000000 101.510000  7.940000 101.660000 ;
      RECT  3.000000 101.510000  7.940000 101.660000 ;
      RECT  3.000000 101.660000  7.795000 101.810000 ;
      RECT  3.000000 101.660000  7.795000 101.810000 ;
      RECT  3.000000 101.810000  7.645000 101.960000 ;
      RECT  3.000000 101.810000  7.645000 101.960000 ;
      RECT  3.000000 101.960000  7.495000 102.110000 ;
      RECT  3.000000 101.960000  7.495000 102.110000 ;
      RECT  3.000000 102.110000  7.345000 102.260000 ;
      RECT  3.000000 102.110000  7.345000 102.260000 ;
      RECT  3.000000 102.260000  7.190000 102.410000 ;
      RECT  3.000000 102.260000  7.190000 102.410000 ;
      RECT  3.000000 102.410000  7.045000 102.560000 ;
      RECT  3.000000 102.410000  7.045000 102.560000 ;
      RECT  3.000000 102.560000  6.895000 102.710000 ;
      RECT  3.000000 102.560000  6.895000 102.710000 ;
      RECT  3.000000 102.710000  6.745000 102.860000 ;
      RECT  3.000000 102.710000  6.745000 102.860000 ;
      RECT  3.000000 102.860000  6.595000 103.010000 ;
      RECT  3.000000 102.860000  6.595000 103.010000 ;
      RECT  3.000000 103.010000  6.440000 103.160000 ;
      RECT  3.000000 103.010000  6.440000 103.160000 ;
      RECT  3.000000 103.160000  6.420000 103.185000 ;
      RECT  3.000000 103.160000  6.420000 103.185000 ;
      RECT  3.000000 122.355000  6.105000 122.505000 ;
      RECT  3.000000 122.355000  6.105000 122.505000 ;
      RECT  3.000000 122.505000  6.255000 122.655000 ;
      RECT  3.000000 122.505000  6.255000 122.655000 ;
      RECT  3.000000 122.655000  6.400000 122.805000 ;
      RECT  3.000000 122.655000  6.400000 122.805000 ;
      RECT  3.000000 122.805000  6.555000 122.955000 ;
      RECT  3.000000 122.805000  6.555000 122.955000 ;
      RECT  3.000000 122.955000  6.705000 123.105000 ;
      RECT  3.000000 122.955000  6.705000 123.105000 ;
      RECT  3.000000 123.105000  6.850000 123.255000 ;
      RECT  3.000000 123.105000  6.850000 123.255000 ;
      RECT  3.000000 123.255000  7.005000 123.405000 ;
      RECT  3.000000 123.255000  7.005000 123.405000 ;
      RECT  3.000000 123.405000  7.150000 123.555000 ;
      RECT  3.000000 123.405000  7.150000 123.555000 ;
      RECT  3.000000 123.555000  7.305000 123.705000 ;
      RECT  3.000000 123.555000  7.305000 123.705000 ;
      RECT  3.000000 123.705000  7.455000 123.855000 ;
      RECT  3.000000 123.705000  7.455000 123.855000 ;
      RECT  3.000000 123.855000  7.600000 124.005000 ;
      RECT  3.000000 123.855000  7.600000 124.005000 ;
      RECT  3.000000 124.005000  7.755000 124.155000 ;
      RECT  3.000000 124.005000  7.755000 124.155000 ;
      RECT  3.000000 124.155000  7.900000 124.305000 ;
      RECT  3.000000 124.155000  7.900000 124.305000 ;
      RECT  3.000000 124.305000  8.055000 124.455000 ;
      RECT  3.000000 124.305000  8.055000 124.455000 ;
      RECT  3.000000 124.455000  8.205000 124.605000 ;
      RECT  3.000000 124.455000  8.205000 124.605000 ;
      RECT  3.000000 124.605000  8.355000 124.650000 ;
      RECT  3.000000 124.605000  8.355000 124.650000 ;
      RECT  3.000000 124.650000 77.000000 172.385000 ;
      RECT  4.455000  73.310000 75.330000  91.880000 ;
      RECT  4.670000   3.000000 75.330000  73.310000 ;
      RECT  4.670000  91.880000 75.330000  98.400000 ;
      RECT  4.670000 172.385000 75.330000 197.000000 ;
      RECT  9.880000 121.400000 12.460000 121.650000 ;
      RECT 12.800000 104.315000 80.000000 121.550000 ;
      RECT 12.900000  95.400000 80.000000 121.650000 ;
      RECT 15.900000 101.210000 77.000000 124.650000 ;
      RECT 75.325000   4.640000 78.330000   7.885000 ;
      RECT 75.325000   7.885000 80.000000   8.485000 ;
      RECT 75.325000   8.485000 78.330000  13.935000 ;
      RECT 75.325000  13.935000 80.000000  14.535000 ;
      RECT 75.325000  14.535000 78.635000  18.785000 ;
      RECT 75.325000  18.785000 80.000000  19.385000 ;
      RECT 75.325000  19.385000 78.330000  24.835000 ;
      RECT 75.325000  24.835000 80.000000  25.435000 ;
      RECT 75.325000  25.435000 78.330000  30.885000 ;
      RECT 75.325000  30.885000 80.000000  31.485000 ;
      RECT 75.325000  31.485000 78.330000  35.735000 ;
      RECT 75.325000  35.735000 80.000000  36.335000 ;
      RECT 75.325000  36.335000 78.330000  40.585000 ;
      RECT 75.325000  40.585000 80.000000  41.185000 ;
      RECT 75.325000  41.185000 78.330000  46.635000 ;
      RECT 75.325000  46.635000 80.000000  47.335000 ;
      RECT 75.325000  47.335000 78.330000  57.135000 ;
      RECT 75.325000  57.135000 80.000000  57.835000 ;
      RECT 75.325000  57.835000 78.330000  63.085000 ;
      RECT 75.325000  63.085000 80.000000  63.685000 ;
      RECT 75.325000  63.685000 78.330000  68.935000 ;
      RECT 75.325000  68.935000 80.000000  69.635000 ;
      RECT 75.325000  69.635000 78.330000  94.885000 ;
      RECT 75.325000 175.385000 78.330000 196.995000 ;
      RECT 75.330000 172.380000 80.000000 175.385000 ;
      RECT 76.995000 121.650000 80.000000 172.380000 ;
    LAYER met5 ;
      RECT  0.000000   0.000000 80.000000 106.585000 ;
      RECT  0.000000 118.955000 80.000000 124.670000 ;
      RECT  0.000000 124.670000 31.315000 147.815000 ;
      RECT  0.000000 147.815000 80.000000 200.000000 ;
      RECT  2.000000 106.585000 80.000000 118.955000 ;
      RECT 54.455000 124.670000 80.000000 147.815000 ;
  END
END sky130_fd_io__top_gpiov2
END LIBRARY
