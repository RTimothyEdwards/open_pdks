magic
tech sky130A
magscale 1 2
timestamp 1607710904
<< metal1 >>
rect 15240 14964 17187 15070
rect 15240 9435 15318 14964
rect 17081 9435 17187 14964
rect 15240 7496 17187 9435
rect 15240 5414 15313 7496
rect 17115 5414 17187 7496
rect 4185 -163 10707 -7
rect 15240 -163 17187 5414
rect 4185 -1384 17187 -163
rect 4185 -2184 16387 -1384
tri 16387 -2184 17187 -1384 nw
<< via1 >>
rect 15318 9435 17081 14964
rect 15313 5414 17115 7496
<< metal2 >>
rect 15240 39521 17187 39586
rect 15240 34813 15294 39521
rect 17136 34813 17187 39521
rect 15240 14964 17187 34813
rect 15240 9435 15318 14964
rect 17081 9435 17187 14964
rect 15240 9312 17187 9435
rect -2195 8808 100 8833
rect -2195 7925 -2165 8808
rect -210 7925 100 8808
rect -2195 7903 100 7925
rect 14940 8809 17228 8840
rect 14940 7939 15154 8809
rect 16192 7939 17228 8809
rect 14940 7910 17228 7939
rect 15240 7496 17187 7560
rect 15240 5644 15313 7496
rect 17115 5644 17187 7496
rect 15240 4807 15278 5644
rect 17134 4807 17187 5644
rect 15240 4678 17187 4807
<< via2 >>
rect 15294 34813 17136 39521
rect -2165 7925 -210 8808
rect 15154 7939 16192 8809
rect 15278 5414 15313 5644
rect 15313 5414 17115 5644
rect 17115 5414 17134 5644
rect 15278 4807 17134 5414
<< metal3 >>
rect 15240 39521 17187 39586
rect 15240 34813 15294 39521
rect 17136 34813 17187 39521
rect 15240 34743 17187 34813
rect -2195 8808 -179 8833
rect -2195 8807 -2165 8808
rect -2195 7924 -2166 8807
rect -210 7925 -179 8808
rect -211 7924 -179 7925
rect -2195 7903 -179 7924
rect 15121 8809 17228 8840
rect 15121 7939 15154 8809
rect 17192 7939 17228 8809
rect 15121 7910 17228 7939
rect 15240 5644 17187 5683
rect 15240 4807 15278 5644
rect 17134 4807 17187 5644
rect 15240 4753 17187 4807
rect 5228 2263 7341 2269
rect 5228 1400 5234 2263
rect 7335 1400 7341 2263
rect 5228 1394 7341 1400
rect 7705 2261 9818 2267
rect 7705 1398 7711 2261
rect 9812 1398 9818 2261
rect 7705 1392 9818 1398
<< via3 >>
rect 15294 34813 17136 39521
rect -2166 7925 -2165 8807
rect -2165 7925 -211 8807
rect -2166 7924 -211 7925
rect 15154 7939 16192 8809
rect 16192 7939 17192 8809
rect 15278 4807 17134 5644
rect 5234 1400 7335 2263
rect 7711 1398 9812 2261
<< metal4 >>
rect 14957 39521 17187 39586
rect 14957 34813 15294 39521
rect 17136 34813 17187 39521
rect 14957 34743 17187 34813
rect -2195 8807 14 8833
rect -2195 7924 -2166 8807
rect -211 7924 14 8807
rect -2195 7903 14 7924
rect 14940 8809 17228 8840
rect 14940 7939 15154 8809
rect 17192 7939 17228 8809
rect 14940 7910 17228 7939
rect 14987 5644 17187 5683
rect 14987 4807 15278 5644
rect 17134 4807 17187 5644
rect 14987 4753 17187 4807
rect 5228 2263 7341 2269
rect 5228 1400 5234 2263
rect 7335 1400 7341 2263
rect 5228 1394 7341 1400
rect 7705 2261 9818 2267
rect 7705 1398 7711 2261
rect 9812 1398 9818 2261
rect 7705 1392 9818 1398
<< properties >>
string FIXED_BBOX 0 -7 15000 39593
<< end >>
