VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__signal_5_sym_hv_local_5term
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__signal_5_sym_hv_local_5term ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.955 BY 12.120 ;
  PIN GATE
    ANTENNAGATEAREA 3.400000 ;
    PORT
      LAYER li1 ;
        RECT 3.310 8.925 4.635 9.335 ;
      LAYER mcon ;
        RECT 3.625 9.065 3.795 9.235 ;
        RECT 3.985 9.065 4.155 9.235 ;
      LAYER met1 ;
        RECT 3.515 8.955 4.260 11.795 ;
    END
  END GATE
  PIN NWELLRING
    ANTENNADIFFAREA 24.296999 ;
    PORT
      LAYER nwell ;
        RECT 0.000 10.760 7.955 12.120 ;
        RECT 0.000 1.360 1.360 10.760 ;
        RECT 6.595 1.360 7.955 10.760 ;
        RECT 0.000 0.000 7.955 1.360 ;
      LAYER li1 ;
        RECT 0.330 11.090 7.625 11.790 ;
        RECT 0.330 1.030 1.030 11.090 ;
        RECT 6.925 1.030 7.625 11.090 ;
        RECT 0.330 0.330 7.625 1.030 ;
      LAYER mcon ;
        RECT 1.535 11.355 1.705 11.525 ;
        RECT 1.895 11.355 2.065 11.525 ;
        RECT 2.255 11.355 2.425 11.525 ;
        RECT 2.615 11.355 2.785 11.525 ;
        RECT 2.975 11.355 3.145 11.525 ;
        RECT 4.795 11.355 4.965 11.525 ;
        RECT 5.155 11.355 5.325 11.525 ;
        RECT 5.515 11.355 5.685 11.525 ;
        RECT 5.875 11.355 6.045 11.525 ;
        RECT 6.235 11.355 6.405 11.525 ;
        RECT 0.595 10.005 0.765 10.175 ;
        RECT 0.595 9.645 0.765 9.815 ;
        RECT 0.595 9.285 0.765 9.455 ;
        RECT 0.595 8.925 0.765 9.095 ;
        RECT 0.595 8.565 0.765 8.735 ;
        RECT 0.595 8.205 0.765 8.375 ;
        RECT 0.595 7.845 0.765 8.015 ;
        RECT 0.595 7.485 0.765 7.655 ;
        RECT 0.595 7.125 0.765 7.295 ;
        RECT 0.595 6.765 0.765 6.935 ;
        RECT 0.595 6.405 0.765 6.575 ;
        RECT 0.595 6.045 0.765 6.215 ;
        RECT 0.595 5.685 0.765 5.855 ;
        RECT 0.595 5.325 0.765 5.495 ;
        RECT 0.595 4.965 0.765 5.135 ;
        RECT 0.595 4.605 0.765 4.775 ;
        RECT 0.595 4.245 0.765 4.415 ;
        RECT 0.595 3.885 0.765 4.055 ;
        RECT 0.595 3.525 0.765 3.695 ;
        RECT 0.595 3.165 0.765 3.335 ;
        RECT 0.595 2.805 0.765 2.975 ;
        RECT 0.595 2.445 0.765 2.615 ;
        RECT 0.595 2.085 0.765 2.255 ;
        RECT 0.595 1.725 0.765 1.895 ;
        RECT 0.595 1.365 0.765 1.535 ;
        RECT 7.190 10.005 7.360 10.175 ;
        RECT 7.190 9.645 7.360 9.815 ;
        RECT 7.190 9.285 7.360 9.455 ;
        RECT 7.190 8.925 7.360 9.095 ;
        RECT 7.190 8.565 7.360 8.735 ;
        RECT 7.190 8.205 7.360 8.375 ;
        RECT 7.190 7.845 7.360 8.015 ;
        RECT 7.190 7.485 7.360 7.655 ;
        RECT 7.190 7.125 7.360 7.295 ;
        RECT 7.190 6.765 7.360 6.935 ;
        RECT 7.190 6.405 7.360 6.575 ;
        RECT 7.190 6.045 7.360 6.215 ;
        RECT 7.190 5.685 7.360 5.855 ;
        RECT 7.190 5.325 7.360 5.495 ;
        RECT 7.190 4.965 7.360 5.135 ;
        RECT 7.190 4.605 7.360 4.775 ;
        RECT 7.190 4.245 7.360 4.415 ;
        RECT 7.190 3.885 7.360 4.055 ;
        RECT 7.190 3.525 7.360 3.695 ;
        RECT 7.190 3.165 7.360 3.335 ;
        RECT 7.190 2.805 7.360 2.975 ;
        RECT 7.190 2.445 7.360 2.615 ;
        RECT 7.190 2.085 7.360 2.255 ;
        RECT 7.190 1.725 7.360 1.895 ;
        RECT 7.190 1.365 7.360 1.535 ;
        RECT 5.590 0.540 5.760 0.710 ;
        RECT 5.950 0.540 6.120 0.710 ;
        RECT 6.310 0.540 6.480 0.710 ;
      LAYER met1 ;
        POLYGON 1.040 11.790 1.040 11.080 0.330 11.080 ;
        RECT 1.040 11.090 3.345 11.790 ;
        RECT 4.430 11.090 6.915 11.790 ;
        RECT 1.040 11.080 1.430 11.090 ;
        POLYGON 1.430 11.090 1.440 11.090 1.430 11.080 ;
        POLYGON 6.445 11.090 6.455 11.090 6.455 11.080 ;
        RECT 6.455 11.080 6.915 11.090 ;
        POLYGON 6.915 11.790 7.625 11.080 6.915 11.080 ;
        RECT 0.330 0.345 1.030 11.080 ;
        POLYGON 1.030 11.080 1.430 11.080 1.030 10.680 ;
        POLYGON 6.455 11.080 6.855 11.080 6.855 10.680 ;
        RECT 6.855 10.680 7.625 11.080 ;
        POLYGON 6.855 10.680 6.915 10.680 6.915 10.620 ;
        RECT 6.915 10.620 7.625 10.680 ;
        POLYGON 6.915 10.620 6.925 10.620 6.925 10.610 ;
        POLYGON 6.925 1.510 6.925 1.030 6.445 1.030 ;
        RECT 6.925 1.040 7.625 10.620 ;
        RECT 6.925 1.030 6.930 1.040 ;
        RECT 5.350 0.345 6.930 1.030 ;
        POLYGON 6.930 1.040 7.625 1.040 6.930 0.345 ;
        RECT 0.330 0.330 1.015 0.345 ;
        RECT 5.350 0.330 6.915 0.345 ;
        POLYGON 6.915 0.345 6.930 0.345 6.915 0.330 ;
    END
  END NWELLRING
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 2.965 3.360 3.505 8.755 ;
      LAYER mcon ;
        RECT 3.105 7.745 3.275 7.915 ;
        RECT 3.105 7.385 3.275 7.555 ;
        RECT 3.105 7.025 3.275 7.195 ;
        RECT 3.105 6.665 3.275 6.835 ;
        RECT 3.105 6.305 3.275 6.475 ;
        RECT 3.105 5.945 3.275 6.115 ;
        RECT 3.105 5.585 3.275 5.755 ;
        RECT 3.105 5.225 3.275 5.395 ;
        RECT 3.105 4.865 3.275 5.035 ;
        RECT 3.105 4.505 3.275 4.675 ;
        RECT 3.105 4.145 3.275 4.315 ;
        RECT 3.105 3.785 3.275 3.955 ;
      LAYER met1 ;
        RECT 2.860 0.330 3.860 8.545 ;
    END
  END VGND
  PIN NBODY
    ANTENNADIFFAREA 13.550600 ;
    PORT
      LAYER pwell ;
        RECT 1.660 1.660 6.295 10.460 ;
      LAYER li1 ;
        RECT 1.790 9.620 6.165 10.330 ;
        RECT 1.790 2.490 2.490 9.620 ;
        RECT 5.465 2.490 6.165 9.620 ;
        RECT 1.790 1.790 6.165 2.490 ;
      LAYER mcon ;
        RECT 2.270 9.845 2.440 10.015 ;
        RECT 2.630 9.845 2.800 10.015 ;
        RECT 2.990 9.845 3.160 10.015 ;
        RECT 4.640 9.845 4.810 10.015 ;
        RECT 5.000 9.845 5.170 10.015 ;
        RECT 5.360 9.845 5.530 10.015 ;
        RECT 1.975 8.845 2.145 9.015 ;
        RECT 1.975 8.485 2.145 8.655 ;
        RECT 1.975 8.125 2.145 8.295 ;
        RECT 1.975 7.765 2.145 7.935 ;
        RECT 1.975 7.405 2.145 7.575 ;
        RECT 1.975 7.045 2.145 7.215 ;
        RECT 1.975 6.685 2.145 6.855 ;
        RECT 1.975 6.325 2.145 6.495 ;
        RECT 1.975 5.965 2.145 6.135 ;
        RECT 1.975 5.605 2.145 5.775 ;
        RECT 1.975 5.245 2.145 5.415 ;
        RECT 1.975 4.885 2.145 5.055 ;
        RECT 1.975 4.525 2.145 4.695 ;
        RECT 1.975 4.165 2.145 4.335 ;
        RECT 1.975 3.805 2.145 3.975 ;
        RECT 1.975 3.445 2.145 3.615 ;
        RECT 1.975 3.085 2.145 3.255 ;
        RECT 1.975 2.725 2.145 2.895 ;
        RECT 1.975 2.365 2.145 2.535 ;
        RECT 5.730 8.845 5.900 9.015 ;
        RECT 5.730 8.485 5.900 8.655 ;
        RECT 5.730 8.125 5.900 8.295 ;
        RECT 5.730 7.765 5.900 7.935 ;
        RECT 5.730 7.405 5.900 7.575 ;
        RECT 5.730 7.045 5.900 7.215 ;
        RECT 5.730 6.685 5.900 6.855 ;
        RECT 5.730 6.325 5.900 6.495 ;
        RECT 5.730 5.965 5.900 6.135 ;
        RECT 5.730 5.605 5.900 5.775 ;
        RECT 5.730 5.245 5.900 5.415 ;
        RECT 5.730 4.885 5.900 5.055 ;
        RECT 5.730 4.525 5.900 4.695 ;
        RECT 5.730 4.165 5.900 4.335 ;
        RECT 5.730 3.805 5.900 3.975 ;
        RECT 5.730 3.445 5.900 3.615 ;
        RECT 5.730 3.085 5.900 3.255 ;
        RECT 5.730 2.725 5.900 2.895 ;
        RECT 5.730 2.365 5.900 2.535 ;
        RECT 1.975 2.005 2.145 2.175 ;
        RECT 5.730 2.005 5.900 2.175 ;
      LAYER met1 ;
        POLYGON 2.120 10.330 2.120 10.000 1.790 10.000 ;
        RECT 2.120 10.000 3.345 10.330 ;
        RECT 1.790 9.505 3.345 10.000 ;
        RECT 4.430 10.000 5.835 10.330 ;
        POLYGON 5.835 10.330 6.165 10.000 5.835 10.000 ;
        RECT 4.430 9.505 6.165 10.000 ;
        RECT 1.790 0.345 2.680 9.505 ;
        POLYGON 2.680 9.505 3.055 9.505 2.680 9.130 ;
        POLYGON 5.060 9.505 5.435 9.505 5.435 9.130 ;
        RECT 5.435 9.130 6.165 9.505 ;
        POLYGON 5.435 9.130 5.465 9.130 5.465 9.100 ;
        RECT 5.465 1.790 6.165 9.130 ;
        RECT 1.790 0.330 2.665 0.345 ;
    END
  END NBODY
  PIN IN
    ANTENNADIFFAREA 3.807000 ;
    PORT
      LAYER li1 ;
        RECT 4.440 3.360 4.980 8.755 ;
      LAYER mcon ;
        RECT 4.575 7.745 4.745 7.915 ;
        RECT 4.575 7.385 4.745 7.555 ;
        RECT 4.575 7.025 4.745 7.195 ;
        RECT 4.575 6.665 4.745 6.835 ;
        RECT 4.575 6.305 4.745 6.475 ;
        RECT 4.575 5.945 4.745 6.115 ;
        RECT 4.575 5.585 4.745 5.755 ;
        RECT 4.575 5.225 4.745 5.395 ;
        RECT 4.575 4.865 4.745 5.035 ;
        RECT 4.575 4.505 4.745 4.675 ;
        RECT 4.575 4.145 4.745 4.315 ;
        RECT 4.575 3.785 4.745 3.955 ;
      LAYER met1 ;
        RECT 4.155 0.330 5.155 8.760 ;
    END
  END IN
  OBS
      LAYER met1 ;
        RECT 1.015 0.330 1.030 0.345 ;
        RECT 2.665 0.330 2.680 0.345 ;
  END
END sky130_fd_io__signal_5_sym_hv_local_5term
END LIBRARY

