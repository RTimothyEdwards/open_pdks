magic
tech sky130A
magscale 1 2
timestamp 1602984771
<< error_p >>
rect 8153 2168 8261 2177
rect 7939 1954 8153 1963
rect 2476 1096 2484 1250
rect 2628 1096 2644 1250
rect 3252 1110 3258 1516
rect 4266 1332 4424 1342
rect 4114 1258 4546 1268
rect 4266 1248 4424 1258
rect 5694 1058 6154 1464
rect 7230 1054 7690 1460
rect 1942 770 1972 812
rect 1942 698 1972 740
rect 7899 190 7979 193
<< dnwell >>
rect 7661 2168 8153 2177
rect 890 206 5190 2104
rect 6796 279 8153 2168
rect 6796 270 7899 279
<< nwell >>
rect 7661 2262 8247 2271
rect 790 1890 5284 2198
rect 790 428 1098 1890
rect 4976 428 5284 1890
rect 790 120 5284 428
rect 6702 1963 8247 2262
rect 6702 1954 7899 1963
rect 6702 492 7010 1954
rect 7939 501 8247 1963
rect 7661 492 8247 501
rect 6702 193 8247 492
rect 6702 184 7899 193
<< nmos >>
rect 3302 1110 3432 1516
rect 4266 1258 4424 1332
<< nsonos >>
rect 1652 1082 1810 1488
rect 1942 1082 2072 1488
rect 3100 1110 3258 1516
rect 4266 1108 4424 1214
rect 5852 1058 6010 1464
rect 7388 1054 7546 1460
rect 1942 740 1972 770
<< ndiff >>
rect 1512 1082 1652 1488
rect 1810 1082 1942 1488
rect 2072 1082 2226 1488
rect 2942 1110 3100 1516
rect 3258 1110 3302 1516
rect 3432 1110 3586 1516
rect 4114 1258 4266 1332
rect 4424 1258 4546 1332
rect 4108 1108 4266 1214
rect 4424 1108 4540 1214
rect 5694 1058 5852 1464
rect 6010 1058 6154 1464
rect 7230 1054 7388 1460
rect 7546 1054 7690 1460
rect 1852 740 1942 770
rect 1972 740 2068 770
<< psubdiff >>
rect 2476 1250 2636 1280
rect 2476 1066 2636 1096
<< psubdiffcont >>
rect 2476 1096 2636 1250
<< poly >>
rect 1652 1488 1810 1598
rect 1942 1488 2072 1606
rect 3100 1516 3258 1626
rect 3302 1516 3432 1634
rect 5852 1464 6010 1574
rect 4266 1332 4424 1358
rect 4266 1214 4424 1258
rect 1652 972 1810 1082
rect 1942 968 2072 1082
rect 3100 1000 3258 1110
rect 3302 996 3432 1110
rect 4266 998 4424 1108
rect 7388 1460 7546 1570
rect 1942 770 1972 968
rect 5852 948 6010 1058
rect 7388 944 7546 1054
rect 1942 682 1972 740
<< locali >>
rect 2476 1250 2636 1280
rect 2476 1066 2636 1096
<< labels >>
flabel comment s -94 846 -88 846 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Tunnel_(Tunm)
flabel comment s 1670 2280 1670 2280 0 FreeSans 560 0 0 0 Use_cif_see_SONOS
flabel comment s -72 658 -72 658 0 FreeSans 560 0 0 0 tunm.1
flabel comment s -92 510 -92 516 0 FreeSans 560 0 0 0 tunm.2
flabel comment s -114 326 -114 328 0 FreeSans 560 0 0 0 tunm.3
flabel comment s -116 178 -116 178 0 FreeSans 560 0 0 0 tunm.4
flabel comment s -120 38 -120 38 0 FreeSans 560 0 0 0 tunm.5
flabel comment s 5920 756 5920 756 0 FreeSans 560 0 0 0 tunm.6a
flabel comment s 1952 564 1952 564 0 FreeSans 560 0 0 0 tunm.7
flabel comment s 1954 868 1954 868 0 FreeSans 560 0 0 0 Incorrect
flabel comment s -134 -80 -134 -80 0 FreeSans 560 0 0 0 tunm.8
flabel comment s 3538 2298 3538 2298 0 FreeSans 560 0 0 0 Use_cif_see_COREID_for_tunm.8
flabel comment s 7405 668 7405 668 0 FreeSans 560 0 0 0 tunm.8
<< properties >>
string FIXED_BBOX 785 110 6460 2201
<< end >>
