magic
tech sky130seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
rect 650 2394 710 51210
tri 650 2369 710 2394 nw
<< end >>
