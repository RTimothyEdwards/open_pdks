magic
tech sky130A
magscale 1 2
timestamp 1605993265
<< properties >>
string LEFclass PAD AREAIO
string FIXED_BBOX 0 0 1000 39593
string GDS_FILE /home/xrex/usr/devel/pdks/sky130A/libs.tech/openlane/custom_cells/gds/sky130_ef_io__disconnect_slice_5um.gds
string GDS_END 226
string GDS_START 158
<< end >>
