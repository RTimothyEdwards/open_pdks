magic
tech sky130A
magscale 1 2
timestamp 1602985534
<< error_p >>
rect -44 786 32 1648
rect 2312 938 2458 1798
rect 3994 922 4884 1732
rect 1875 -865 2215 -769
rect 4369 -1187 4763 -377
<< dnwell >>
rect 1657 -1285 2421 -659
rect 3943 -1187 4763 -377
<< nwell >>
rect -215 1648 54 1883
rect -136 786 -44 1648
rect 1340 938 2204 1798
rect 2312 938 3198 1798
rect 3994 922 4884 1732
rect 1519 -769 2555 -430
rect 1519 -1073 1875 -769
rect 2215 -1073 2555 -769
rect 1519 -1401 2555 -1073
rect 3815 -1323 4891 -229
rect 5269 -1147 5959 -433
<< nsubdiff >>
rect -168 1822 9 1844
rect -168 1707 -136 1822
rect -26 1707 9 1822
rect -168 1684 9 1707
rect 1414 1673 1596 1697
rect 1414 1558 1449 1673
rect 1559 1558 1596 1673
rect 1414 1534 1596 1558
rect 2864 1627 3042 1651
rect 2864 1512 2901 1627
rect 3011 1512 3042 1627
rect 2864 1489 3042 1512
rect 3864 -314 4047 -289
rect 3864 -429 3907 -314
rect 4017 -429 4047 -314
rect 3864 -458 4047 -429
rect 1578 -505 1765 -482
rect 1578 -620 1603 -505
rect 1713 -620 1765 -505
rect 1578 -647 1765 -620
rect 5727 -492 5902 -470
rect 5727 -607 5758 -492
rect 5868 -607 5902 -492
rect 5727 -631 5902 -607
<< nsubdiffcont >>
rect -136 1707 -26 1822
rect 1449 1558 1559 1673
rect 2901 1512 3011 1627
rect 3907 -429 4017 -314
rect 1603 -620 1713 -505
rect 5758 -607 5868 -492
<< locali >>
rect -161 1707 -136 1822
rect -26 1707 9 1822
rect -161 1706 9 1707
rect 1419 1558 1449 1673
rect 1559 1558 1588 1673
rect 2872 1627 3039 1628
rect 2872 1512 2901 1627
rect 3011 1512 3039 1627
rect 3867 -429 3907 -314
rect 4017 -429 4069 -314
rect 5707 -492 5916 -491
rect 1558 -620 1603 -505
rect 1713 -620 1756 -505
rect 5707 -607 5758 -492
rect 5868 -607 5916 -492
rect 5707 -608 5916 -607
<< labels >>
flabel comment s 50 -918 50 -918 0 FreeSans 560 0 0 0 (not_implemented)
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Nwell
flabel comment s 2350 802 2350 802 0 FreeSans 560 0 0 0 nwell.2
flabel comment s -78 572 -78 572 0 FreeSans 560 0 0 0 nwell.1
flabel comment s 64 -1108 64 -1108 0 FreeSans 560 0 0 0 nwell.2b
flabel comment s 4340 762 4340 762 0 FreeSans 560 0 0 0 nwell.4
flabel comment s 58 -1252 58 -1252 0 FreeSans 560 0 0 0 nwell.5a
flabel comment s 34 -1390 34 -1390 0 FreeSans 560 0 0 0 nwell.5b
flabel comment s 1983 -1497 1983 -1497 0 FreeSans 560 0 0 0 nwell.6
flabel comment s 4397 -1443 4397 -1443 0 FreeSans 560 0 0 0 nwell.7
<< end >>
