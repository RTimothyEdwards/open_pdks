magic
tech s8seal_ring
magscale 1 2
timestamp 1584562315
<< type81_52 >>
rect 0 20320 20320 51210
rect 0 0 51200 20320
use sr_polygon00028  sr_polygon00028_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 650 2369 710 51210
use sr_polygon00024  sr_polygon00024_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 530 2319 590 51210
use sr_polygon00020  sr_polygon00020_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 410 2269 470 51210
use sr_polygon00016  sr_polygon00016_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 290 2219 350 51210
use sr_polygon00032  sr_polygon00032_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 0 2099 1000 51210
use sr_polygon00031  sr_polygon00031_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 650 650 51200 2394
use sr_polygon00027  sr_polygon00027_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 530 530 51200 2344
use sr_polygon00023  sr_polygon00023_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 410 410 51200 2294
use sr_polygon00019  sr_polygon00019_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 290 290 51200 2244
use nikon_sealring_shape  nikon_sealring_shape_0
timestamp 1584558468
transform 1 0 200 0 1 200
box 0 0 800 800
use sr_polygon00036  sr_polygon00036_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 0 0 1200 51210
use sr_polygon00015  sr_polygon00015_0
timestamp 1584558468
transform 1 0 0 0 1 0
box 0 0 2099 2099
use sr_polygon00035  sr_polygon00035_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 0 0 51200 2514
use sr_polygon00039  sr_polygon00039_0
timestamp 1584558827
transform 1 0 0 0 1 0
box 0 0 51200 2597
use sr_polygon00011  sr_polygon00011_0
timestamp 1584558468
transform 1 0 0 0 1 0
box -30480 -30480 30480 30480
<< end >>
