magic
tech sky130A
magscale 1 2
timestamp 1636577591
<< metal1 >>
rect 15240 14964 17187 15070
rect 15240 9668 15318 14964
rect 17081 9668 17187 14964
rect 15240 5414 15313 9668
rect 17115 5414 17187 9668
rect 5101 -7 5685 83
rect 4185 -163 11313 -7
rect 15240 -163 17187 5414
rect 4185 -1384 17187 -163
rect 4185 -2184 16387 -1384
tri 16387 -2184 17187 -1384 nw
<< via1 >>
rect 15318 9668 17081 14964
rect 15313 5414 17115 9668
<< metal2 >>
rect 15240 39521 17187 39586
rect 15240 34813 15294 39521
rect 17136 34813 17187 39521
rect 15240 14964 17187 34813
rect 15240 9668 15318 14964
rect 17081 9668 17187 14964
rect 15240 5644 15313 9668
rect 17115 5644 17187 9668
rect 15240 4807 15278 5644
rect 17134 4807 17187 5644
rect 15240 4678 17187 4807
<< via2 >>
rect 15294 34813 17136 39521
rect 15278 5414 15313 5644
rect 15313 5414 17115 5644
rect 17115 5414 17134 5644
rect 15278 4807 17134 5414
<< metal3 >>
rect 15240 39521 17187 39586
rect 15240 34813 15294 39521
rect 17136 34813 17187 39521
rect 15240 34743 17187 34813
rect 15240 5644 17187 5683
rect 15240 4807 15278 5644
rect 17134 4807 17187 5644
rect 15240 4753 17187 4807
<< via3 >>
rect 15294 34813 17136 39521
rect 15278 4807 17134 5644
<< metal4 >>
rect 14957 39521 17187 39586
rect 14957 34813 15294 39521
rect 17136 34813 17187 39521
rect 14957 34743 17187 34813
rect 14987 5644 17187 5683
rect 14987 4807 15278 5644
rect 17134 4807 17187 5644
rect 14987 4753 17187 4807
<< properties >>
string FIXED_BBOX 0 -7 15000 39593
<< end >>
