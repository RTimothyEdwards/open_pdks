magic
tech sky130A
magscale 1 2
timestamp 1584473789
<< metal2 >>
rect 99 -407 4879 -259
rect 5179 -407 5579 -181
rect 10078 -407 14858 -259
<< metal3 >>
rect 99 -407 4879 -16
rect 5179 -407 7379 -259
rect 7578 -407 9778 -89
rect 10078 -407 14858 -16
<< metal4 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 0 13600 254 18593
rect 14746 13600 15000 18593
rect 0 12410 254 13300
rect 14746 12410 15000 13300
rect 0 11240 254 12130
rect 14746 11240 15000 12130
rect 0 10874 254 10940
rect 14746 10874 15000 10940
rect 0 10218 100 10814
rect 14746 10218 14846 10814
rect 0 9922 254 10158
rect 14746 9922 15000 10158
rect 0 9266 116 9862
rect 14746 9266 14862 9862
rect 0 9140 254 9206
rect 14746 9140 15000 9206
rect 0 7910 254 8840
rect 14746 7910 15000 8840
rect 0 6940 254 7630
rect 14746 6940 15000 7630
rect 0 5970 254 6660
rect 14746 5970 15000 6660
rect 0 4760 254 5690
rect 14746 4760 15000 5690
rect 0 3550 254 4480
rect 14746 3550 15000 4480
rect 0 2580 254 3270
rect 14746 2580 15000 3270
rect 0 1370 254 2300
rect 14746 1370 15000 2300
rect 0 6 254 1090
rect 14746 6 15000 1090
rect 14934 5 15000 6
rect 0 0 254 5
rect 14746 0 15000 5
<< metal5 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 7329 27458 7594 28780
rect 0 13600 254 18590
rect 14746 13600 15000 18590
rect 0 12430 254 13280
rect 14746 12430 15000 13280
rect 0 11260 254 12110
rect 14746 11260 15000 12110
rect 0 9140 254 10940
rect 14746 9140 15000 10940
rect 0 7930 254 8820
rect 14746 7930 15000 8820
rect 0 6960 254 7610
rect 14746 6960 15000 7610
rect 0 5990 254 6640
rect 14746 5990 15000 6640
rect 0 4780 254 5670
rect 14746 4780 15000 5670
rect 0 3570 254 4460
rect 14746 3570 15000 4460
rect 0 2600 254 3250
rect 14746 2600 15000 3250
rect 0 1390 254 2280
rect 14746 1390 15000 2280
rect 0 20 254 1070
rect 14746 20 15000 1070
use sky130_fd_io__overlay_vssio_hvc  sky130_fd_io__overlay_vssio_hvc_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1584046481
transform 1 0 0 0 1 -407
box 0 407 15000 40000
use sky130_fd_io__top_ground_hvc_wpad  sky130_fd_io__top_ground_hvc_wpad_2 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1584046481
transform 1 0 0 0 1 -407
box 0 0 15000 40000
<< labels >>
flabel metal5 s 7329 27458 7594 28780 0 FreeSans 2000 0 0 0 vssio
port 12 nsew
flabel metal4 s 127 37914 127 37914 3 FreeSans 520 0 0 0 vssio
port 12 nsew
flabel metal4 s 14873 37914 14873 37914 3 FreeSans 520 180 0 0 vssio
port 12 nsew
flabel metal2 s 10078 -407 14858 -259 2 FreeSans 2000 90 0 0 drn_hvc
port 2 nsew
flabel metal2 s 99 -407 4879 -259 2 FreeSans 2000 90 0 0 src_bdy_hvc
port 4 nsew
flabel metal3 s 7578 -407 9778 -89 0 FreeSans 2000 0 0 0 drn_hvc
port 2 nsew
flabel metal3 s 99 -407 4879 -16 0 FreeSans 2000 0 0 0 vssio
port 12 nsew
flabel metal3 s 10078 -407 14858 -16 0 FreeSans 2000 0 0 0 vssio
port 12 nsew
flabel metal3 s 5179 -407 7379 -259 2 FreeSans 2000 90 0 0 src_bdy_hvc
port 4 nsew
flabel metal5 s 14746 9140 15000 10940 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal5 s 14807 2600 15000 3250 3 FreeSans 520 180 0 0 vdda
port 6 nsew
flabel metal5 s 14746 7930 15000 8820 3 FreeSans 520 180 0 0 vssd
port 13 nsew
flabel metal5 s 14746 11260 15000 12110 3 FreeSans 520 180 0 0 vssio_q
port 14 nsew
flabel metal5 s 14746 4780 15000 5670 3 FreeSans 520 180 0 0 vssio
port 12 nsew
flabel metal5 s 14746 5990 15000 6640 3 FreeSans 520 180 0 0 vswitch
port 7 nsew
flabel metal5 s 14746 6961 15000 7610 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal5 s 14746 1390 15000 2280 3 FreeSans 520 180 0 0 vccd
port 11 nsew
flabel metal5 s 14746 12430 15000 13280 3 FreeSans 520 180 0 0 vddio_q
port 8 nsew
flabel metal5 s 14746 13600 15000 18590 3 FreeSans 520 180 0 0 vddio
port 10 nsew
flabel metal5 s 14746 20 15000 1070 3 FreeSans 520 180 0 0 vcchib
port 9 nsew
flabel metal5 s 14746 3570 15000 4460 3 FreeSans 520 180 0 0 vddio
port 10 nsew
flabel metal5 s 0 13600 254 18590 3 FreeSans 520 0 0 0 vddio
port 10 nsew
flabel metal5 s 0 7930 254 8820 3 FreeSans 520 0 0 0 vssd
port 13 nsew
flabel metal5 s 0 11260 254 12110 3 FreeSans 520 0 0 0 vssio_q
port 14 nsew
flabel metal5 s 0 5990 254 6640 3 FreeSans 520 0 0 0 vswitch
port 7 nsew
flabel metal5 s 0 4780 254 5670 3 FreeSans 520 0 0 0 vssio
port 12 nsew
flabel metal5 s 0 2600 193 3250 3 FreeSans 520 0 0 0 vdda
port 6 nsew
flabel metal5 s 0 3570 254 4460 3 FreeSans 520 0 0 0 vddio
port 10 nsew
flabel metal5 s 0 1390 254 2280 3 FreeSans 520 0 0 0 vccd
port 11 nsew
flabel metal5 s 0 12430 254 13280 3 FreeSans 520 0 0 0 vddio_q
port 8 nsew
flabel metal5 s 0 9140 254 10940 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal5 s 0 6961 254 7610 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal5 s 0 20 254 1070 3 FreeSans 520 0 0 0 vcchib
port 9 nsew
flabel metal4 s 14746 7910 15000 8840 3 FreeSans 520 180 0 0 vssd
port 13 nsew
flabel metal4 s 14807 2580 15000 3270 3 FreeSans 520 180 0 0 vdda
port 6 nsew
flabel metal4 s 14746 11240 15000 12130 3 FreeSans 520 180 0 0 vssio_q
port 14 nsew
flabel metal4 s 14746 4760 15000 5690 3 FreeSans 520 180 0 0 vssio
port 12 nsew
flabel metal4 s 14746 5970 15000 6660 3 FreeSans 520 180 0 0 vswitch
port 7 nsew
flabel metal4 s 14746 9922 15000 10158 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 14746 10874 15000 10940 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 14746 0 15000 1090 3 FreeSans 520 180 0 0 vcchib
port 9 nsew
flabel metal4 s 14746 3550 15000 4480 3 FreeSans 520 180 0 0 vddio
port 10 nsew
flabel metal4 s 14746 9140 15000 9206 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 14746 6940 15000 7630 3 FreeSans 520 180 0 0 vssa
port 5 nsew
flabel metal4 s 14746 12410 15000 13300 3 FreeSans 520 180 0 0 vddio_q
port 8 nsew
flabel metal4 s 14746 1370 15000 2300 3 FreeSans 520 180 0 0 vccd
port 11 nsew
flabel metal4 s 14746 9266 15000 9862 3 FreeSans 520 180 0 0 amuxbus_b
port 1 nsew
flabel metal4 s 14746 34750 15000 39593 3 FreeSans 520 180 0 0 vssio
port 12 nsew
flabel metal4 s 14746 10218 15000 10814 3 FreeSans 520 180 0 0 amuxbus_a
port 0 nsew
flabel metal4 s 14746 13600 15000 18593 3 FreeSans 520 180 0 0 vddio
port 10 nsew
flabel metal4 s 0 34750 254 39593 3 FreeSans 520 0 0 0 vssio
port 12 nsew
flabel metal4 s 0 3550 254 4480 3 FreeSans 520 0 0 0 vddio
port 10 nsew
flabel metal4 s 0 12410 254 13300 3 FreeSans 520 0 0 0 vddio_q
port 8 nsew
flabel metal4 s 0 13600 254 18593 3 FreeSans 520 0 0 0 vddio
port 10 nsew
flabel metal4 s 0 1370 254 2300 3 FreeSans 520 0 0 0 vccd
port 11 nsew
flabel metal4 s 0 9140 254 9206 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 5970 254 6660 3 FreeSans 520 0 0 0 vswitch
port 7 nsew
flabel metal4 s 0 0 254 1090 3 FreeSans 520 0 0 0 vcchib
port 9 nsew
flabel metal4 s 0 9922 254 10158 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 11240 254 12130 3 FreeSans 520 0 0 0 vssio_q
port 14 nsew
flabel metal4 s 0 4760 254 5690 3 FreeSans 520 0 0 0 vssio
port 12 nsew
flabel metal4 s 0 2580 193 3270 3 FreeSans 520 0 0 0 vdda
port 6 nsew
flabel metal4 s 0 10218 254 10814 3 FreeSans 520 0 0 0 amuxbus_a
port 0 nsew
flabel metal4 s 0 10874 254 10940 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 6940 254 7630 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal4 s 0 7910 254 8840 3 FreeSans 520 0 0 0 vssd
port 13 nsew
flabel metal4 s 0 9266 254 9862 3 FreeSans 520 0 0 0 amuxbus_b
port 1 nsew
<< properties >>
string LEFclass PAD GROUND
string FIXED_BBOX 0 0 15000 39593
<< end >>
