magic
tech sky130A
magscale 1 2
timestamp 1602597384
<< error_s >>
rect 1668 39147 1734 39163
rect 2691 37377 2692 37401
rect 2772 37377 2773 37401
rect 3245 37377 3246 37401
rect 3326 37377 3327 37401
rect 3799 37377 3800 37401
rect 3880 37377 3881 37401
rect 4353 37377 4354 37401
rect 4434 37377 4435 37401
rect 4907 37377 4908 37401
rect 4988 37377 4989 37401
rect 5461 37377 5462 37401
rect 5542 37377 5543 37401
rect 6015 37377 6016 37401
rect 6096 37377 6097 37401
rect 6569 37377 6570 37401
rect 6650 37377 6651 37401
rect 7123 37377 7124 37401
rect 7204 37377 7205 37401
rect 7677 37377 7678 37401
rect 7758 37377 7759 37401
rect 8231 37377 8232 37401
rect 8312 37377 8313 37401
rect 8785 37377 8786 37401
rect 8866 37377 8867 37401
rect 9339 37377 9340 37401
rect 9420 37377 9421 37401
rect 9893 37377 9894 37401
rect 9974 37377 9975 37401
rect 10447 37377 10448 37401
rect 10528 37377 10529 37401
rect 11001 37377 11002 37401
rect 11082 37377 11083 37401
rect 11555 37377 11556 37401
rect 11636 37377 11637 37401
rect 12109 37377 12110 37401
rect 12190 37377 12191 37401
rect 12663 37377 12664 37401
rect 12744 37377 12745 37401
rect 13217 37377 13218 37401
rect 13298 37377 13299 37401
rect 2715 37353 2749 37365
rect 3269 37353 3303 37365
rect 3823 37353 3857 37365
rect 4377 37353 4411 37365
rect 4931 37353 4965 37365
rect 5485 37353 5519 37365
rect 6039 37353 6073 37365
rect 6593 37353 6627 37365
rect 7147 37353 7181 37365
rect 7701 37353 7735 37365
rect 8255 37353 8289 37365
rect 8809 37353 8843 37365
rect 9363 37353 9397 37365
rect 9917 37353 9951 37365
rect 10471 37353 10505 37365
rect 11025 37353 11059 37365
rect 11579 37353 11613 37365
rect 12133 37353 12167 37365
rect 12687 37353 12721 37365
rect 13241 37353 13275 37365
rect 3245 35377 3246 35401
rect 3326 35377 3327 35401
rect 3799 35377 3800 35401
rect 3880 35377 3881 35401
rect 4353 35377 4354 35401
rect 4434 35377 4435 35401
rect 4907 35377 4908 35401
rect 4988 35377 4989 35401
rect 5461 35377 5462 35401
rect 5542 35377 5543 35401
rect 6015 35377 6016 35401
rect 6096 35377 6097 35401
rect 6569 35377 6570 35401
rect 6650 35377 6651 35401
rect 7123 35377 7124 35401
rect 7204 35377 7205 35401
rect 7677 35377 7678 35401
rect 7758 35377 7759 35401
rect 8231 35377 8232 35401
rect 8312 35377 8313 35401
rect 8785 35377 8786 35401
rect 8866 35377 8867 35401
rect 9339 35377 9340 35401
rect 9420 35377 9421 35401
rect 9893 35377 9894 35401
rect 9974 35377 9975 35401
rect 10447 35377 10448 35401
rect 10528 35377 10529 35401
rect 11001 35377 11002 35401
rect 11082 35377 11083 35401
rect 11555 35377 11556 35401
rect 11636 35377 11637 35401
rect 12109 35377 12110 35401
rect 12190 35377 12191 35401
rect 12663 35377 12664 35401
rect 12744 35377 12745 35401
rect 13217 35377 13218 35401
rect 13298 35377 13299 35401
rect 3269 35353 3303 35365
rect 3823 35353 3857 35365
rect 4377 35353 4411 35365
rect 4931 35353 4965 35365
rect 5485 35353 5519 35365
rect 6039 35353 6073 35365
rect 6593 35353 6627 35365
rect 7147 35353 7181 35365
rect 7701 35353 7735 35365
rect 8255 35353 8289 35365
rect 8809 35353 8843 35365
rect 9363 35353 9397 35365
rect 9917 35353 9951 35365
rect 10471 35353 10505 35365
rect 11025 35353 11059 35365
rect 11579 35353 11613 35365
rect 12133 35353 12167 35365
rect 12687 35353 12721 35365
rect 13241 35353 13275 35365
rect 3185 33377 3186 33401
rect 3266 33377 3267 33401
rect 4021 33377 4022 33401
rect 4102 33377 4103 33401
rect 4857 33377 4858 33401
rect 4938 33377 4939 33401
rect 5693 33377 5694 33401
rect 5774 33377 5775 33401
rect 6529 33377 6530 33401
rect 6610 33377 6611 33401
rect 7365 33377 7366 33401
rect 7446 33377 7447 33401
rect 8201 33377 8202 33401
rect 8282 33377 8283 33401
rect 9037 33377 9038 33401
rect 9118 33377 9119 33401
rect 9873 33377 9874 33401
rect 9954 33377 9955 33401
rect 10709 33377 10710 33401
rect 10790 33377 10791 33401
rect 11545 33377 11546 33401
rect 11626 33377 11627 33401
rect 12381 33377 12382 33401
rect 12462 33377 12463 33401
rect 13217 33377 13218 33401
rect 13298 33377 13299 33401
rect 3209 33353 3243 33365
rect 4045 33353 4079 33365
rect 4881 33353 4915 33365
rect 5717 33353 5751 33365
rect 6553 33353 6587 33365
rect 7389 33353 7423 33365
rect 8225 33353 8259 33365
rect 9061 33353 9095 33365
rect 9897 33353 9931 33365
rect 10733 33353 10767 33365
rect 11569 33353 11603 33365
rect 12405 33353 12439 33365
rect 13241 33353 13275 33365
rect 3185 31377 3186 31401
rect 3266 31377 3267 31401
rect 4021 31377 4022 31401
rect 4102 31377 4103 31401
rect 4857 31377 4858 31401
rect 4938 31377 4939 31401
rect 5693 31377 5694 31401
rect 5774 31377 5775 31401
rect 6529 31377 6530 31401
rect 6610 31377 6611 31401
rect 7365 31377 7366 31401
rect 7446 31377 7447 31401
rect 8201 31377 8202 31401
rect 8282 31377 8283 31401
rect 9037 31377 9038 31401
rect 9118 31377 9119 31401
rect 9873 31377 9874 31401
rect 9954 31377 9955 31401
rect 10709 31377 10710 31401
rect 10790 31377 10791 31401
rect 11545 31377 11546 31401
rect 11626 31377 11627 31401
rect 12381 31377 12382 31401
rect 12462 31377 12463 31401
rect 13217 31377 13218 31401
rect 13298 31377 13299 31401
rect 3209 31353 3243 31365
rect 4045 31353 4079 31365
rect 4881 31353 4915 31365
rect 5717 31353 5751 31365
rect 6553 31353 6587 31365
rect 7389 31353 7423 31365
rect 8225 31353 8259 31365
rect 9061 31353 9095 31365
rect 9897 31353 9931 31365
rect 10733 31353 10767 31365
rect 11569 31353 11603 31365
rect 12405 31353 12439 31365
rect 13241 31353 13275 31365
rect 3185 29377 3186 29401
rect 3266 29377 3267 29401
rect 4021 29377 4022 29401
rect 4102 29377 4103 29401
rect 4857 29377 4858 29401
rect 4938 29377 4939 29401
rect 5693 29377 5694 29401
rect 5774 29377 5775 29401
rect 6529 29377 6530 29401
rect 6610 29377 6611 29401
rect 7365 29377 7366 29401
rect 7446 29377 7447 29401
rect 8201 29377 8202 29401
rect 8282 29377 8283 29401
rect 9037 29377 9038 29401
rect 9118 29377 9119 29401
rect 9873 29377 9874 29401
rect 9954 29377 9955 29401
rect 10709 29377 10710 29401
rect 10790 29377 10791 29401
rect 11545 29377 11546 29401
rect 11626 29377 11627 29401
rect 12381 29377 12382 29401
rect 12462 29377 12463 29401
rect 13217 29377 13218 29401
rect 13298 29377 13299 29401
rect 3209 29353 3243 29365
rect 4045 29353 4079 29365
rect 4881 29353 4915 29365
rect 5717 29353 5751 29365
rect 6553 29353 6587 29365
rect 7389 29353 7423 29365
rect 8225 29353 8259 29365
rect 9061 29353 9095 29365
rect 9897 29353 9931 29365
rect 10733 29353 10767 29365
rect 11569 29353 11603 29365
rect 12405 29353 12439 29365
rect 13241 29353 13275 29365
rect 4857 27377 4858 27401
rect 4938 27377 4939 27401
rect 5693 27377 5694 27401
rect 5774 27377 5775 27401
rect 6529 27377 6530 27401
rect 6610 27377 6611 27401
rect 7365 27377 7366 27401
rect 7446 27377 7447 27401
rect 8201 27377 8202 27401
rect 8282 27377 8283 27401
rect 9037 27377 9038 27401
rect 9118 27377 9119 27401
rect 9873 27377 9874 27401
rect 9954 27377 9955 27401
rect 10709 27377 10710 27401
rect 10790 27377 10791 27401
rect 11545 27377 11546 27401
rect 11626 27377 11627 27401
rect 12381 27377 12382 27401
rect 12462 27377 12463 27401
rect 13217 27377 13218 27401
rect 13298 27377 13299 27401
rect 4881 27353 4915 27365
rect 5717 27353 5751 27365
rect 6553 27353 6587 27365
rect 7389 27353 7423 27365
rect 8225 27353 8259 27365
rect 9061 27353 9095 27365
rect 9897 27353 9931 27365
rect 10733 27353 10767 27365
rect 11569 27353 11603 27365
rect 12405 27353 12439 27365
rect 13241 27353 13275 27365
rect 4857 25756 4858 25780
rect 4938 25756 4939 25780
rect 5693 25756 5694 25780
rect 5774 25756 5775 25780
rect 6529 25756 6530 25780
rect 6610 25756 6611 25780
rect 7365 25756 7366 25780
rect 7446 25756 7447 25780
rect 8201 25756 8202 25780
rect 8282 25756 8283 25780
rect 9037 25756 9038 25780
rect 9118 25756 9119 25780
rect 9873 25756 9874 25780
rect 9954 25756 9955 25780
rect 10709 25756 10710 25780
rect 10790 25756 10791 25780
rect 11545 25756 11546 25780
rect 11626 25756 11627 25780
rect 12381 25756 12382 25780
rect 12462 25756 12463 25780
rect 13217 25756 13218 25780
rect 13298 25756 13299 25780
rect 4881 25732 4915 25744
rect 5717 25732 5751 25744
rect 6553 25732 6587 25744
rect 7389 25732 7423 25744
rect 8225 25732 8259 25744
rect 9061 25732 9095 25744
rect 9897 25732 9931 25744
rect 10733 25732 10767 25744
rect 11569 25732 11603 25744
rect 12405 25732 12439 25744
rect 13241 25732 13275 25744
rect 2691 13377 2692 13401
rect 2772 13377 2773 13401
rect 3245 13377 3246 13401
rect 3326 13377 3327 13401
rect 3799 13377 3800 13401
rect 3880 13377 3881 13401
rect 4353 13377 4354 13401
rect 4434 13377 4435 13401
rect 4907 13377 4908 13401
rect 4988 13377 4989 13401
rect 5461 13377 5462 13401
rect 5542 13377 5543 13401
rect 6015 13377 6016 13401
rect 6096 13377 6097 13401
rect 6569 13377 6570 13401
rect 6650 13377 6651 13401
rect 7123 13377 7124 13401
rect 7204 13377 7205 13401
rect 7677 13377 7678 13401
rect 7758 13377 7759 13401
rect 8231 13377 8232 13401
rect 8312 13377 8313 13401
rect 8785 13377 8786 13401
rect 8866 13377 8867 13401
rect 9339 13377 9340 13401
rect 9420 13377 9421 13401
rect 9893 13377 9894 13401
rect 9974 13377 9975 13401
rect 10447 13377 10448 13401
rect 10528 13377 10529 13401
rect 11001 13377 11002 13401
rect 11082 13377 11083 13401
rect 11555 13377 11556 13401
rect 11636 13377 11637 13401
rect 12109 13377 12110 13401
rect 12190 13377 12191 13401
rect 12663 13377 12664 13401
rect 12744 13377 12745 13401
rect 13217 13377 13218 13401
rect 13298 13377 13299 13401
rect 2715 13353 2749 13365
rect 3269 13353 3303 13365
rect 3823 13353 3857 13365
rect 4377 13353 4411 13365
rect 4931 13353 4965 13365
rect 5485 13353 5519 13365
rect 6039 13353 6073 13365
rect 6593 13353 6627 13365
rect 7147 13353 7181 13365
rect 7701 13353 7735 13365
rect 8255 13353 8289 13365
rect 8809 13353 8843 13365
rect 9363 13353 9397 13365
rect 9917 13353 9951 13365
rect 10471 13353 10505 13365
rect 11025 13353 11059 13365
rect 11579 13353 11613 13365
rect 12133 13353 12167 13365
rect 12687 13353 12721 13365
rect 13241 13353 13275 13365
rect 2691 11377 2692 11401
rect 2772 11377 2773 11401
rect 3245 11377 3246 11401
rect 3326 11377 3327 11401
rect 3799 11377 3800 11401
rect 3880 11377 3881 11401
rect 4353 11377 4354 11401
rect 4434 11377 4435 11401
rect 4907 11377 4908 11401
rect 4988 11377 4989 11401
rect 5461 11377 5462 11401
rect 5542 11377 5543 11401
rect 6015 11377 6016 11401
rect 6096 11377 6097 11401
rect 6569 11377 6570 11401
rect 6650 11377 6651 11401
rect 7123 11377 7124 11401
rect 7204 11377 7205 11401
rect 7677 11377 7678 11401
rect 7758 11377 7759 11401
rect 8231 11377 8232 11401
rect 8312 11377 8313 11401
rect 8785 11377 8786 11401
rect 8866 11377 8867 11401
rect 9339 11377 9340 11401
rect 9420 11377 9421 11401
rect 9893 11377 9894 11401
rect 9974 11377 9975 11401
rect 10447 11377 10448 11401
rect 10528 11377 10529 11401
rect 11001 11377 11002 11401
rect 11082 11377 11083 11401
rect 11555 11377 11556 11401
rect 11636 11377 11637 11401
rect 12109 11377 12110 11401
rect 12190 11377 12191 11401
rect 12663 11377 12664 11401
rect 12744 11377 12745 11401
rect 13217 11377 13218 11401
rect 13298 11377 13299 11401
rect 2715 11353 2749 11365
rect 3269 11353 3303 11365
rect 3823 11353 3857 11365
rect 4377 11353 4411 11365
rect 4931 11353 4965 11365
rect 5485 11353 5519 11365
rect 6039 11353 6073 11365
rect 6593 11353 6627 11365
rect 7147 11353 7181 11365
rect 7701 11353 7735 11365
rect 8255 11353 8289 11365
rect 8809 11353 8843 11365
rect 9363 11353 9397 11365
rect 9917 11353 9951 11365
rect 10471 11353 10505 11365
rect 11025 11353 11059 11365
rect 11579 11353 11613 11365
rect 12133 11353 12167 11365
rect 12687 11353 12721 11365
rect 13241 11353 13275 11365
rect 2691 9377 2692 9401
rect 2772 9377 2773 9401
rect 3245 9377 3246 9401
rect 3326 9377 3327 9401
rect 3799 9377 3800 9401
rect 3880 9377 3881 9401
rect 4353 9377 4354 9401
rect 4434 9377 4435 9401
rect 4907 9377 4908 9401
rect 4988 9377 4989 9401
rect 5461 9377 5462 9401
rect 5542 9377 5543 9401
rect 6015 9377 6016 9401
rect 6096 9377 6097 9401
rect 6569 9377 6570 9401
rect 6650 9377 6651 9401
rect 7123 9377 7124 9401
rect 7204 9377 7205 9401
rect 7677 9377 7678 9401
rect 7758 9377 7759 9401
rect 8231 9377 8232 9401
rect 8312 9377 8313 9401
rect 8785 9377 8786 9401
rect 8866 9377 8867 9401
rect 9339 9377 9340 9401
rect 9420 9377 9421 9401
rect 9893 9377 9894 9401
rect 9974 9377 9975 9401
rect 10447 9377 10448 9401
rect 10528 9377 10529 9401
rect 11001 9377 11002 9401
rect 11082 9377 11083 9401
rect 11555 9377 11556 9401
rect 11636 9377 11637 9401
rect 12109 9377 12110 9401
rect 12190 9377 12191 9401
rect 12663 9377 12664 9401
rect 12744 9377 12745 9401
rect 13217 9377 13218 9401
rect 13298 9377 13299 9401
rect 2715 9353 2749 9365
rect 3269 9353 3303 9365
rect 3823 9353 3857 9365
rect 4377 9353 4411 9365
rect 4931 9353 4965 9365
rect 5485 9353 5519 9365
rect 6039 9353 6073 9365
rect 6593 9353 6627 9365
rect 7147 9353 7181 9365
rect 7701 9353 7735 9365
rect 8255 9353 8289 9365
rect 8809 9353 8843 9365
rect 9363 9353 9397 9365
rect 9917 9353 9951 9365
rect 10471 9353 10505 9365
rect 11025 9353 11059 9365
rect 11579 9353 11613 9365
rect 12133 9353 12167 9365
rect 12687 9353 12721 9365
rect 13241 9353 13275 9365
rect 2691 7377 2692 7401
rect 2772 7377 2773 7401
rect 3245 7377 3246 7401
rect 3326 7377 3327 7401
rect 3799 7377 3800 7401
rect 3880 7377 3881 7401
rect 4353 7377 4354 7401
rect 4434 7377 4435 7401
rect 4907 7377 4908 7401
rect 4988 7377 4989 7401
rect 5461 7377 5462 7401
rect 5542 7377 5543 7401
rect 6015 7377 6016 7401
rect 6096 7377 6097 7401
rect 6569 7377 6570 7401
rect 6650 7377 6651 7401
rect 7123 7377 7124 7401
rect 7204 7377 7205 7401
rect 7677 7377 7678 7401
rect 7758 7377 7759 7401
rect 8231 7377 8232 7401
rect 8312 7377 8313 7401
rect 8785 7377 8786 7401
rect 8866 7377 8867 7401
rect 9339 7377 9340 7401
rect 9420 7377 9421 7401
rect 9893 7377 9894 7401
rect 9974 7377 9975 7401
rect 10447 7377 10448 7401
rect 10528 7377 10529 7401
rect 11001 7377 11002 7401
rect 11082 7377 11083 7401
rect 11555 7377 11556 7401
rect 11636 7377 11637 7401
rect 12109 7377 12110 7401
rect 12190 7377 12191 7401
rect 12663 7377 12664 7401
rect 12744 7377 12745 7401
rect 13217 7377 13218 7401
rect 13298 7377 13299 7401
rect 2715 7353 2749 7365
rect 3269 7353 3303 7365
rect 3823 7353 3857 7365
rect 4377 7353 4411 7365
rect 4931 7353 4965 7365
rect 5485 7353 5519 7365
rect 6039 7353 6073 7365
rect 6593 7353 6627 7365
rect 7147 7353 7181 7365
rect 7701 7353 7735 7365
rect 8255 7353 8289 7365
rect 8809 7353 8843 7365
rect 9363 7353 9397 7365
rect 9917 7353 9951 7365
rect 10471 7353 10505 7365
rect 11025 7353 11059 7365
rect 11579 7353 11613 7365
rect 12133 7353 12167 7365
rect 12687 7353 12721 7365
rect 13241 7353 13275 7365
rect 2691 5377 2692 5401
rect 2772 5377 2773 5401
rect 3245 5377 3246 5401
rect 3326 5377 3327 5401
rect 3799 5377 3800 5401
rect 3880 5377 3881 5401
rect 4353 5377 4354 5401
rect 4434 5377 4435 5401
rect 4907 5377 4908 5401
rect 4988 5377 4989 5401
rect 5461 5377 5462 5401
rect 5542 5377 5543 5401
rect 6015 5377 6016 5401
rect 6096 5377 6097 5401
rect 6569 5377 6570 5401
rect 6650 5377 6651 5401
rect 7123 5377 7124 5401
rect 7204 5377 7205 5401
rect 7677 5377 7678 5401
rect 7758 5377 7759 5401
rect 8231 5377 8232 5401
rect 8312 5377 8313 5401
rect 8785 5377 8786 5401
rect 8866 5377 8867 5401
rect 9339 5377 9340 5401
rect 9420 5377 9421 5401
rect 9893 5377 9894 5401
rect 9974 5377 9975 5401
rect 10447 5377 10448 5401
rect 10528 5377 10529 5401
rect 11001 5377 11002 5401
rect 11082 5377 11083 5401
rect 11555 5377 11556 5401
rect 11636 5377 11637 5401
rect 12109 5377 12110 5401
rect 12190 5377 12191 5401
rect 12663 5377 12664 5401
rect 12744 5377 12745 5401
rect 13217 5377 13218 5401
rect 13298 5377 13299 5401
rect 2715 5353 2749 5365
rect 3269 5353 3303 5365
rect 3823 5353 3857 5365
rect 4377 5353 4411 5365
rect 4931 5353 4965 5365
rect 5485 5353 5519 5365
rect 6039 5353 6073 5365
rect 6593 5353 6627 5365
rect 7147 5353 7181 5365
rect 7701 5353 7735 5365
rect 8255 5353 8289 5365
rect 8809 5353 8843 5365
rect 9363 5353 9397 5365
rect 9917 5353 9951 5365
rect 10471 5353 10505 5365
rect 11025 5353 11059 5365
rect 11579 5353 11613 5365
rect 12133 5353 12167 5365
rect 12687 5353 12721 5365
rect 13241 5353 13275 5365
rect 48 3833 114 3849
rect 7279 3663 7365 3699
rect 3525 469 3825 3469
rect 3968 3414 4206 3438
rect 3968 548 3969 3414
rect 3944 525 3969 548
rect 4206 525 4230 3414
rect 3944 524 4230 525
rect 3968 500 3992 524
rect 4349 469 4649 3469
rect 4792 3414 5030 3438
rect 4792 548 4793 3414
rect 4768 525 4793 548
rect 5030 525 5054 3414
rect 4768 524 5054 525
rect 4792 500 4816 524
rect 5173 469 5473 3469
rect 5616 3414 5854 3438
rect 5616 548 5617 3414
rect 5592 525 5617 548
rect 5854 525 5878 3414
rect 5592 524 5878 525
rect 5616 500 5640 524
rect 5997 469 6297 3469
rect 6440 3414 6678 3438
rect 6440 548 6441 3414
rect 6416 525 6441 548
rect 6678 525 6702 3414
rect 6416 524 6702 525
rect 6440 500 6464 524
rect 6821 469 7121 3469
rect 7279 275 7315 3663
rect 7329 275 7365 3663
rect 7523 469 7823 3469
rect 7966 3414 8204 3438
rect 7966 548 7967 3414
rect 7942 525 7967 548
rect 8204 525 8228 3414
rect 7942 524 8228 525
rect 7966 500 7990 524
rect 8347 469 8647 3469
rect 8790 3414 9028 3438
rect 8790 548 8791 3414
rect 8766 525 8791 548
rect 9028 525 9052 3414
rect 8766 524 9052 525
rect 8790 500 8814 524
rect 9171 469 9471 3469
rect 9614 3414 9852 3438
rect 9614 548 9615 3414
rect 9590 525 9615 548
rect 9852 525 9876 3414
rect 9590 524 9876 525
rect 9614 500 9638 524
rect 9995 469 10295 3469
rect 10438 3414 10676 3438
rect 10438 548 10439 3414
rect 10414 525 10439 548
rect 10676 525 10700 3414
rect 10414 524 10700 525
rect 10438 500 10462 524
rect 10819 469 11119 3469
rect 7279 239 7365 275
<< metal1 >>
rect 6867 95 7067 195
rect 5242 -7 5540 74
<< metal2 >>
rect 100 0 4099 287
rect 6888 -7 8888 58
rect 10953 -7 14940 715
<< metal3 >>
rect 98 339 4900 862
rect 100 0 4900 339
rect 5200 -7 7374 918
rect 7676 -7 9850 918
rect 10151 -7 14940 862
<< metal4 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 0 13600 254 18593
rect 14746 13600 15000 18593
rect 0 12410 254 13300
rect 14746 12410 15000 13300
rect 0 11240 254 12130
rect 14746 11240 15000 12130
rect 0 10874 254 10940
rect 14746 10874 15000 10940
rect 0 10218 100 10814
rect 14746 10218 14846 10814
rect 0 9922 254 10158
rect 14746 9922 15000 10158
rect 0 9266 116 9862
rect 14746 9266 14862 9862
rect 0 9140 254 9206
rect 14746 9140 15000 9206
rect 0 7910 254 8840
rect 14746 7910 15000 8840
rect 0 6940 254 7630
rect 14746 6940 15000 7630
rect 0 5970 254 6660
rect 14746 5970 15000 6660
rect 0 4760 254 5690
rect 14746 4760 15000 5690
rect 0 3550 254 4480
rect 14746 3550 15000 4480
rect 0 2580 254 3270
rect 14746 2580 15000 3270
rect 0 1370 254 2300
rect 14746 1370 15000 2300
rect 0 0 254 1090
rect 14746 0 15000 1090
<< metal5 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 6339 32546 10468 33417
rect 0 13600 254 18590
rect 14746 13600 15000 18590
rect 0 12430 254 13280
rect 14746 12430 15000 13280
rect 0 11260 254 12110
rect 14746 11260 15000 12110
rect 0 9140 254 10940
rect 14746 9140 15000 10940
rect 0 7930 254 8820
rect 14746 7930 15000 8820
rect 0 6960 254 7610
rect 14746 6960 15000 7610
rect 0 5990 254 6640
rect 14746 5990 15000 6640
rect 0 4780 254 5670
rect 14746 4780 15000 5670
rect 0 3570 254 4460
rect 14746 3570 15000 4460
rect 0 2600 254 3250
rect 14746 2600 15000 3250
rect 0 1390 254 2280
rect 14746 1390 15000 2280
rect 0 20 254 1070
rect 14746 20 15000 1070
use sky130_fd_io__top_ground_lvc_wpad  sky130_fd_io__top_ground_lvc_wpad_2 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602555073
transform 1 0 0 0 1 -7
box 0 0 15000 39600
use sky130_fd_io__overlay_vssio_lvc  sky130_fd_io__overlay_vssio_lvc_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602555073
transform 1 0 0 0 1 -7
box 0 7 15000 39600
<< labels >>
flabel metal5 s 6339 32546 10468 33417 0 FreeSans 2000 0 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal2 s 100 -7 4099 287 0 FreeSans 2000 0 0 0 SRC_BDY_LVC1
port 4 nsew ground bidirectional
flabel metal2 s 10953 -7 14940 715 0 FreeSans 2000 0 0 0 SRC_BDY_LVC2
port 5 nsew ground bidirectional
flabel metal2 s 6888 -7 8888 58 0 FreeSans 400 0 0 0 BDY2_B2B
port 6 nsew ground bidirectional
flabel metal3 s 7676 -7 9850 918 0 FreeSans 2000 0 0 0 DRN_LVC2
port 3 nsew power bidirectional
flabel metal3 s 5200 -7 7374 918 0 FreeSans 2000 0 0 0 DRN_LVC1
port 2 nsew power bidirectional
flabel metal3 s 10151 -7 14940 862 0 FreeSans 4000 0 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal3 s 100 -7 4900 862 0 FreeSans 2000 0 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal5 s 14746 9140 15000 10940 3 FreeSans 520 180 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal5 s 14807 2600 15000 3250 3 FreeSans 520 180 0 0 VDDA
port 10 nsew power bidirectional
flabel metal5 s 14746 7930 15000 8820 3 FreeSans 520 180 0 0 VSSD
port 17 nsew ground bidirectional
flabel metal5 s 14746 11260 15000 12110 3 FreeSans 520 180 0 0 VSSIO_Q
port 18 nsew ground bidirectional
flabel metal5 s 14746 4780 15000 5670 3 FreeSans 520 180 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal5 s 14746 5990 15000 6640 3 FreeSans 520 180 0 0 VSWITCH
port 11 nsew power bidirectional
flabel metal5 s 14746 6961 15000 7610 3 FreeSans 520 180 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal5 s 14746 1390 15000 2280 3 FreeSans 520 180 0 0 VCCD
port 15 nsew power bidirectional
flabel metal5 s 14746 12430 15000 13280 3 FreeSans 520 180 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal5 s 14746 13600 15000 18590 3 FreeSans 520 180 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal5 s 14746 20 15000 1070 3 FreeSans 520 180 0 0 VCCHIB
port 13 nsew power bidirectional
flabel metal5 s 14746 3570 15000 4460 3 FreeSans 520 180 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal5 s 0 13600 254 18590 3 FreeSans 520 0 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal5 s 0 7930 254 8820 3 FreeSans 520 0 0 0 VSSD
port 17 nsew ground bidirectional
flabel metal5 s 0 11260 254 12110 3 FreeSans 520 0 0 0 VSSIO_Q
port 18 nsew ground bidirectional
flabel metal5 s 0 5990 254 6640 3 FreeSans 520 0 0 0 VSWITCH
port 11 nsew power bidirectional
flabel metal5 s 0 4780 254 5670 3 FreeSans 520 0 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal5 s 0 2600 193 3250 3 FreeSans 520 0 0 0 VDDA
port 10 nsew power bidirectional
flabel metal5 s 0 3570 254 4460 3 FreeSans 520 0 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal5 s 0 1390 254 2280 3 FreeSans 520 0 0 0 VCCD
port 15 nsew power bidirectional
flabel metal5 s 0 12430 254 13280 3 FreeSans 520 0 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal5 s 0 9140 254 10940 3 FreeSans 520 0 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal5 s 0 6961 254 7610 3 FreeSans 520 0 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal5 s 0 20 254 1070 3 FreeSans 520 0 0 0 VCCHIB
port 13 nsew power bidirectional
flabel metal4 s 14746 7910 15000 8840 3 FreeSans 520 180 0 0 VSSD
port 17 nsew ground bidirectional
flabel metal4 s 14807 2580 15000 3270 3 FreeSans 520 180 0 0 VDDA
port 10 nsew power bidirectional
flabel metal4 s 14746 11240 15000 12130 3 FreeSans 520 180 0 0 VSSIO_Q
port 18 nsew ground bidirectional
flabel metal4 s 14746 4760 15000 5690 3 FreeSans 520 180 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal4 s 14746 5970 15000 6660 3 FreeSans 520 180 0 0 VSWITCH
port 11 nsew power bidirectional
flabel metal4 s 14746 9922 15000 10158 3 FreeSans 520 180 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 14746 10874 15000 10940 3 FreeSans 520 180 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 14746 0 15000 1090 3 FreeSans 520 180 0 0 VCCHIB
port 13 nsew power bidirectional
flabel metal4 s 14746 3550 15000 4480 3 FreeSans 520 180 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal4 s 14746 9140 15000 9206 3 FreeSans 520 180 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 14746 6940 15000 7630 3 FreeSans 520 180 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 14746 12410 15000 13300 3 FreeSans 520 180 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal4 s 14746 1370 15000 2300 3 FreeSans 520 180 0 0 VCCD
port 15 nsew power bidirectional
flabel metal4 s 14746 9266 15000 9862 3 FreeSans 520 180 0 0 AMUXBUS_B
port 1 nsew signal bidirectional
flabel metal4 s 14746 34750 15000 39593 3 FreeSans 520 180 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal4 s 14746 10218 15000 10814 3 FreeSans 520 180 0 0 AMUXBUS_A
port 0 nsew signal bidirectional
flabel metal4 s 14746 13600 15000 18593 3 FreeSans 520 180 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal4 s 0 34750 254 39593 3 FreeSans 520 0 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal4 s 0 3550 254 4480 3 FreeSans 520 0 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal4 s 0 12410 254 13300 3 FreeSans 520 0 0 0 VDDIO_Q
port 12 nsew power bidirectional
flabel metal4 s 0 13600 254 18593 3 FreeSans 520 0 0 0 VDDIO
port 14 nsew power bidirectional
flabel metal4 s 0 1370 254 2300 3 FreeSans 520 0 0 0 VCCD
port 15 nsew power bidirectional
flabel metal4 s 0 9140 254 9206 3 FreeSans 520 0 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 0 5970 254 6660 3 FreeSans 520 0 0 0 VSWITCH
port 11 nsew power bidirectional
flabel metal4 s 0 0 254 1090 3 FreeSans 520 0 0 0 VCCHIB
port 13 nsew power bidirectional
flabel metal4 s 0 9922 254 10158 3 FreeSans 520 0 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 0 11240 254 12130 3 FreeSans 520 0 0 0 VSSIO_Q
port 18 nsew ground bidirectional
flabel metal4 s 0 4760 254 5690 3 FreeSans 520 0 0 0 VSSIO
port 16 nsew ground bidirectional
flabel metal4 s 0 2580 193 3270 3 FreeSans 520 0 0 0 VDDA
port 10 nsew power bidirectional
flabel metal4 s 0 10218 254 10814 3 FreeSans 520 0 0 0 AMUXBUS_A
port 0 nsew signal bidirectional
flabel metal4 s 0 10874 254 10940 3 FreeSans 520 0 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 0 6940 254 7630 3 FreeSans 520 0 0 0 VSSA
port 9 nsew ground bidirectional
flabel metal4 s 0 7910 254 8840 3 FreeSans 520 0 0 0 VSSD
port 17 nsew ground bidirectional
flabel metal4 s 0 9266 254 9862 3 FreeSans 520 0 0 0 AMUXBUS_B
port 1 nsew signal bidirectional
<< properties >>
string LEFclass PAD GROUND
string FIXED_BBOX 0 0 15000 39593
<< end >>
