* NGSPICE file created from sky130_ef_io__analog_pad.ext - technology: sky130A

.subckt sky130_fd_io__pad_esd m4_960_20017# m5_1354_20500#
R0 m4_960_20017# m5_1354_20500# sky130_fd_pr__res_generic_m5 w=253 l=0.1
.ends

.subckt sky130_fd_io__com_busses_esd sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__com_bus_hookup_0/VSSD
+ sky130_fd_io__pad_esd_0/m5_1354_20500# sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__pad_esd_0/m4_960_20017#
+ sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_bus_hookup_0/VCCD
Xsky130_fd_io__pad_esd_0 sky130_fd_io__pad_esd_0/m4_960_20017# sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__pad_esd
.ends

.subckt sky130_ef_io__esd_pdiode_11v0_array a_n1540_n5136# a_1132_n5000# a_516_n5000#
+ a_n1332_n5000# a_n716_n5000# a_n100_n5000#
D0 a_n716_n5000# a_n716_n5000# sky130_fd_pr__diode_pw2nd_11v0 pj=1.02e+08 area=5e+13
D1 a_n1332_n5000# a_n1332_n5000# sky130_fd_pr__diode_pw2nd_11v0 pj=1.02e+08 area=5e+13
D2 a_n100_n5000# a_n100_n5000# sky130_fd_pr__diode_pw2nd_11v0 pj=1.02e+08 area=5e+13
D3 a_1132_n5000# a_1132_n5000# sky130_fd_pr__diode_pw2nd_11v0 pj=1.02e+08 area=5e+13
D4 a_516_n5000# a_516_n5000# sky130_fd_pr__diode_pw2nd_11v0 pj=1.02e+08 area=5e+13
.ends

.subckt sky130_ef_io__esd_ndiode_11v0_array a_964_n5000# a_n1164_n5000# a_432_n5000#
+ a_n632_n5000# a_n100_n5000# w_n1396_n5168#
D0 a_432_n5000# w_n1396_n5168# sky130_fd_pr__diode_pd2nw_11v0 pj=1.02e+08 area=5e+13
D1 a_n100_n5000# w_n1396_n5168# sky130_fd_pr__diode_pd2nw_11v0 pj=1.02e+08 area=5e+13
D2 a_n632_n5000# w_n1396_n5168# sky130_fd_pr__diode_pd2nw_11v0 pj=1.02e+08 area=5e+13
D3 a_964_n5000# w_n1396_n5168# sky130_fd_pr__diode_pd2nw_11v0 pj=1.02e+08 area=5e+13
D4 a_n1164_n5000# w_n1396_n5168# sky130_fd_pr__diode_pd2nw_11v0 pj=1.02e+08 area=5e+13
.ends

.subckt sky130_ef_io__esd_pad_and_busses sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
+ m1_2509_27880# sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH
Xsky130_fd_io__com_busses_esd_0 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA
+ m1_2509_27880# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_busses_esd
Xsky130_ef_io__esd_vssio sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ m1_2509_27880# m1_2509_27880# m1_2509_27880# m1_2509_27880# m1_2509_27880# sky130_ef_io__esd_pdiode_11v0_array
Xsky130_ef_io__esd_vddio m1_2509_27880# m1_2509_27880# m1_2509_27880# m1_2509_27880#
+ m1_2509_27880# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO
+ sky130_ef_io__esd_ndiode_11v0_array
.ends

.subckt sky130_ef_io__analog_pad P_CORE VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO
+ VSWITCH VSSIO VDDA VCCD VCCHIB VSSIO_Q P_PAD
Xsky130_ef_io__esd_pad_and_busses_0 VCCD P_CORE P_PAD VSSD VDDIO_Q VSSA AMUXBUS_B
+ AMUXBUS_A VSSIO_Q VDDIO VCCHIB VSSIO VDDA VSWITCH sky130_ef_io__esd_pad_and_busses
.ends

