magic
tech sky130A
magscale 1 2
timestamp 1597519380
<< error_p >>
rect 1249 1260 1333 1268
<< nmos >>
rect 1266 1144 1313 1230
rect 1499 1144 1529 1230
rect 1631 1144 1661 1230
<< ndiff >>
rect 1185 1144 1266 1230
rect 1313 1144 1499 1230
rect 1529 1144 1631 1230
rect 1661 1144 1721 1230
<< poly >>
rect 1233 1347 1349 1357
rect 1233 1260 1249 1347
rect 1333 1260 1349 1347
rect 1233 1250 1349 1260
rect 1481 1302 1547 1312
rect 1481 1268 1497 1302
rect 1531 1268 1547 1302
rect 1481 1258 1547 1268
rect 1621 1302 1675 1318
rect 1621 1268 1631 1302
rect 1665 1268 1675 1302
rect 1266 1230 1313 1250
rect 1499 1230 1529 1258
rect 1621 1252 1675 1268
rect 1631 1230 1661 1252
rect 1932 1214 1998 1224
rect 1932 1180 1948 1214
rect 1982 1180 1998 1214
rect 1932 1170 1998 1180
rect 1266 1100 1313 1144
rect 1499 1114 1529 1144
rect 1631 1114 1661 1144
rect 1837 1127 1903 1137
rect 1837 1093 1853 1127
rect 1887 1093 1903 1127
rect 1837 1083 1903 1093
<< polycont >>
rect 1249 1260 1333 1347
rect 1497 1268 1531 1302
rect 1631 1268 1665 1302
rect 1948 1180 1982 1214
rect 1853 1093 1887 1127
<< locali >>
rect 1193 1260 1249 1347
rect 1333 1260 1393 1347
rect 1441 1268 1497 1302
rect 1531 1268 1631 1302
rect 1665 1268 1716 1302
rect 1892 1180 1948 1214
rect 1982 1180 2042 1214
rect 1797 1093 1853 1127
rect 1887 1093 1947 1127
<< labels >>
flabel comment s -23 575 -17 575 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s -15 1143 -9 1143 0 FreeSans 560 0 0 0 Not_Implemented
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Nitride_Poly_Cut_(npc)
flabel comment s 1626 2208 1626 2208 0 FreeSans 560 0 0 0 Use_cif_see_NPC
flabel comment s -39 354 -39 354 0 FreeSans 560 0 0 0 npc.1
flabel comment s -19 185 -19 185 0 FreeSans 560 0 0 0 npc.2
flabel comment s -19 -60 -19 -60 0 FreeSans 560 0 0 0 npc.3
flabel comment s 1289 907 1289 907 0 FreeSans 560 0 0 0 npc.4
flabel comment s 23 893 23 893 0 FreeSans 560 0 0 0 npc.5
<< end >>
