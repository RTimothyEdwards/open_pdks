* Power pads library (s8 power pads + overlays)
* Includes corner and fill cell subcircuits

.SUBCKT s8iom0_vdda_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vdda_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vddio_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vddio_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vccd_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vccd_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vssa_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vssa_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vssio_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vssio_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vssd_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_vssd_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_corner_pad
+ amuxbus_a amuxbus_b 
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0s8_com_bus_slice
+ amuxbus_a amuxbus_b
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0s8_com_bus_slice_1um
+ amuxbus_a amuxbus_b
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT s8iom0_gpiov2_pad
+ in_h pad_a_noesd_h pad_a_esd_0_h pad_a_esd_1_h
+ pad dm<2> dm<1> dm<0> hld_h_n in inp_dis ib_mode_sel enable_h enable_vdda_h
+ enable_inp_h oe_n tie_hi_esd tie_lo_esd slow vtrip_sel hld_ovr
+ analog_en analog_sel enable_vddio enable_vswitch_h analog_pol out
+ amuxbus_a amuxbus_b vssa vdda vswitch vddio_q vcchib vddio vccd vssio
+ vssd vssio_q
.ENDS
