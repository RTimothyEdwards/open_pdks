magic
tech sky130seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
tri 290 2219 350 2244 se
tri 350 2219 375 2244 sw
tri 290 2134 375 2219 ne
tri 375 2134 460 2219 sw
tri 375 2049 460 2134 ne
tri 460 2049 545 2134 sw
tri 460 1964 545 2049 ne
tri 545 1964 630 2049 sw
tri 545 1879 630 1964 ne
tri 630 1879 715 1964 sw
tri 630 1794 715 1879 ne
tri 715 1794 800 1879 sw
tri 715 1709 800 1794 ne
tri 800 1709 885 1794 sw
tri 800 1624 885 1709 ne
tri 885 1624 970 1709 sw
tri 885 1539 970 1624 ne
tri 970 1539 1055 1624 sw
tri 970 1454 1055 1539 ne
tri 1055 1454 1140 1539 sw
tri 1055 1369 1140 1454 ne
tri 1140 1369 1225 1454 sw
tri 1140 1284 1225 1369 ne
tri 1225 1284 1310 1369 sw
tri 1225 1199 1310 1284 ne
tri 1310 1199 1395 1284 sw
tri 1310 1114 1395 1199 ne
tri 1395 1114 1480 1199 sw
tri 1395 1029 1480 1114 ne
tri 1480 1029 1565 1114 sw
tri 1480 944 1565 1029 ne
tri 1565 944 1650 1029 sw
tri 1565 859 1650 944 ne
tri 1650 859 1735 944 sw
tri 1650 774 1735 859 ne
tri 1735 774 1820 859 sw
tri 1735 689 1820 774 ne
tri 1820 689 1905 774 sw
tri 1820 604 1905 689 ne
tri 1905 604 1990 689 sw
tri 1905 519 1990 604 ne
tri 1990 519 2075 604 sw
tri 1990 434 2075 519 ne
tri 2075 434 2160 519 sw
tri 2075 349 2160 434 ne
tri 2160 350 2244 434 sw
rect 2160 349 51200 350
tri 2160 290 2219 349 ne
rect 2219 290 51200 349
<< end >>
