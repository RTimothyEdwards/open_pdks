magic
tech sky130seal_ring
magscale 1 2
timestamp 1584558827
<< type61_20 >>
rect 0 2514 1000 51210
tri 0 2099 1000 2514 nw
<< end >>
