magic
tech sky130A
timestamp 1607711116
<< metal3 >>
rect 2640 19728 3633 19731
rect 1454 19723 2447 19726
rect 368 19720 1364 19723
rect 368 18362 371 19720
rect 1361 18362 1364 19720
rect 368 18359 1364 18362
rect 1454 17436 1457 19723
rect 2444 17436 2447 19723
rect 2640 17441 2643 19728
rect 3630 17441 3633 19728
rect 2640 17438 3633 17441
rect 1454 17433 2447 17436
rect 3812 9272 4873 9275
rect 3812 6825 3815 9272
rect 4870 6825 4873 9272
rect 3812 6822 4873 6825
rect 2608 2827 3668 2830
rect 2608 2399 2611 2827
rect 3665 2399 3668 2827
rect 2608 2396 3668 2399
rect 3802 2222 4875 2225
rect 3802 1795 3805 2222
rect 4872 1795 4875 2222
rect 3802 1792 4875 1795
<< via3 >>
rect 371 18362 1361 19720
rect 1457 17436 2444 19723
rect 2643 17441 3630 19728
rect 3815 6825 4870 9272
rect 2611 2399 3665 2827
rect 3805 1795 4872 2222
<< metal4 >>
rect 2640 19728 3633 19731
rect 1454 19723 2447 19726
rect 368 19720 1364 19723
rect 368 18362 371 19720
rect 1361 18362 1364 19720
rect 368 18359 1364 18362
rect 1454 17436 1457 19723
rect 2444 17436 2447 19723
rect 2640 17441 2643 19728
rect 3630 17441 3633 19728
rect 2640 17438 3633 17441
rect 1454 17433 2447 17436
rect 3812 9272 4873 9275
rect 3812 6825 3815 9272
rect 4870 6825 4873 9272
rect 3812 6822 4873 6825
rect 2608 2827 3668 2830
rect 2608 2399 2611 2827
rect 3665 2399 3668 2827
rect 2608 2396 3668 2399
rect 3802 2222 4875 2225
rect 3802 1795 3805 2222
rect 4872 1795 4875 2222
rect 3802 1792 4875 1795
<< properties >>
string FIXED_BBOX 0 -203 7500 19796
<< end >>
