magic
tech sky130seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
rect 530 2344 590 51210
tri 530 2319 590 2344 nw
<< end >>
