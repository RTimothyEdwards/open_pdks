* For diodes called as a subcircuit
* (backwards compatible with earlier PDK version)
.subckt sky130_fd_pr__diode_pw2nd N P a=0 p=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=a
.ends
* (corresponds to current PDK)
.subckt sky130_fd_pr__diode_pw2nd_05v5 N P area=0
D0 N P sky130_fd_pr__diode_pw2nd_05v5 area=area
.ends
