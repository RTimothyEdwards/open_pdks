magic
tech sky130A
magscale 1 2
timestamp 1602970101
<< error_p >>
rect 2560 930 2568 1084
rect 2712 930 2728 1084
rect 3332 944 3342 1350
rect 6336 1206 6390 1346
rect 6424 1206 6478 1346
rect 4350 1102 4508 1120
rect 5978 862 5986 1016
rect 6130 862 6146 1016
rect 8238 894 8344 1300
rect 8602 908 8610 1062
rect 8754 908 8770 1062
rect 2504 -782 2512 -628
rect 2656 -782 2672 -628
rect 3278 -768 3286 -362
rect 7904 -422 7912 -268
rect 8056 -422 8072 -268
rect 4294 -610 4452 -592
rect 6524 -652 6578 -500
rect 6592 -652 6646 -500
rect 8014 -714 8025 -703
rect 8137 -714 8148 -703
rect 6162 -1002 6170 -848
rect 6314 -1002 6330 -848
rect 8003 -910 8014 -899
rect 8148 -910 8159 -899
<< nwell >>
rect 1386 708 4858 1660
rect 5790 704 6980 1762
rect 7522 686 8866 1638
rect 7774 -1022 8476 -138
<< pwell >>
rect 1326 -1208 5166 -122
rect 5914 -1224 7104 -166
<< nmos >>
rect 3361 -768 3491 -362
rect 4294 -610 4452 -546
<< pmos >>
rect 3415 944 3545 1350
rect 4350 1102 4508 1166
<< mvvaractor >>
rect 8014 -910 8148 -714
<< pmoslvt >>
rect 1736 916 1894 1322
rect 2026 916 2156 1322
rect 3184 944 3342 1350
rect 4350 942 4508 1048
rect 8238 894 8396 1300
rect 6524 -652 6592 -500
<< pmoshvt >>
rect 8116 894 8196 1300
<< nmoslvt >>
rect 6336 1206 6424 1346
rect 1680 -796 1838 -390
rect 1970 -796 2100 -390
rect 3128 -768 3286 -362
rect 4294 -770 4452 -664
<< ndiff >>
rect 1540 -796 1680 -390
rect 1838 -796 1970 -390
rect 2100 -796 2254 -390
rect 2970 -768 3128 -362
rect 3286 -768 3361 -362
rect 3491 -768 3645 -362
rect 4142 -610 4294 -546
rect 4452 -610 4574 -546
rect 6354 -652 6524 -500
rect 6592 -652 6796 -500
rect 4136 -770 4294 -664
rect 4452 -770 4568 -664
<< pdiff >>
rect 1596 916 1736 1322
rect 1894 916 2026 1322
rect 2156 916 2310 1322
rect 3026 944 3184 1350
rect 3342 944 3415 1350
rect 3545 944 3699 1350
rect 6144 1206 6336 1346
rect 6424 1206 6672 1346
rect 4198 1102 4350 1166
rect 4508 1102 4630 1166
rect 4192 942 4350 1048
rect 4508 942 4624 1048
rect 8018 894 8116 1300
rect 8196 894 8238 1300
rect 8396 894 8438 1300
<< psubdiff >>
rect 2504 -628 2664 -598
rect 2504 -812 2664 -782
rect 6162 -848 6322 -818
rect 6162 -1032 6322 -1002
<< nsubdiff >>
rect 2560 1084 2720 1114
rect 2560 900 2720 930
rect 5978 1016 6138 1046
rect 8602 1062 8762 1092
rect 5978 832 6138 862
rect 8602 878 8762 908
rect 7904 -268 8064 -238
rect 7904 -452 8064 -422
<< mvnsubdiff >>
rect 7932 -910 8014 -714
rect 8148 -910 8230 -714
<< psubdiffcont >>
rect 2504 -782 2664 -628
rect 6162 -1002 6322 -848
<< nsubdiffcont >>
rect 2560 930 2720 1084
rect 5978 862 6138 1016
rect 8602 908 8762 1062
rect 7904 -422 8064 -268
<< poly >>
rect 1736 1322 1894 1432
rect 2026 1322 2156 1440
rect 3184 1350 3342 1460
rect 3415 1350 3545 1468
rect 6336 1346 6424 1452
rect 8116 1300 8196 1408
rect 8238 1300 8396 1410
rect 4350 1166 4508 1192
rect 4350 1048 4508 1102
rect 6336 1086 6424 1206
rect 1736 806 1894 916
rect 2026 802 2156 916
rect 3184 834 3342 944
rect 3415 830 3545 944
rect 4350 832 4508 942
rect 8116 780 8196 894
rect 8238 784 8396 894
rect 1680 -390 1838 -280
rect 1970 -390 2100 -272
rect 3128 -362 3286 -252
rect 3361 -362 3491 -244
rect 6524 -500 6592 -380
rect 4294 -546 4452 -520
rect 4294 -664 4452 -610
rect 1680 -906 1838 -796
rect 1970 -910 2100 -796
rect 3128 -878 3286 -768
rect 3361 -882 3491 -768
rect 6524 -752 6592 -652
rect 8014 -714 8148 -662
rect 4294 -880 4452 -770
rect 8014 -962 8148 -910
<< locali >>
rect 2560 1084 2720 1114
rect 8602 1062 8762 1092
rect 2560 900 2720 930
rect 5978 1016 6138 1046
rect 8602 878 8762 908
rect 5978 832 6138 862
rect 7904 -268 8064 -238
rect 7904 -452 8064 -422
rect 2504 -628 2664 -598
rect 2504 -812 2664 -782
rect 6162 -848 6322 -818
rect 6162 -1032 6322 -1002
<< labels >>
flabel comment s -94 846 -88 846 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Lvtn_(Lvtnm)
flabel comment s -72 658 -72 658 0 FreeSans 560 0 0 0 lvtn.1
flabel comment s -92 510 -92 516 0 FreeSans 560 0 0 0 lvtn.2
flabel comment s 1670 2280 1670 2280 0 FreeSans 560 0 0 0 Use_cif_see_LVTN
flabel comment s 8152 572 8152 572 0 FreeSans 560 0 0 0 lvtn.9
flabel comment s -114 326 -114 328 0 FreeSans 560 0 0 0 lvtn.3b
flabel comment s -120 166 -120 166 0 FreeSans 560 0 0 0 lvtn.13
flabel comment s -140 -12 -140 -12 0 FreeSans 560 0 0 0 lvtn.14
flabel comment s -144 -188 -144 -188 0 FreeSans 560 0 0 0 lvtn.12
flabel comment s 3342 587 3342 587 0 FreeSans 560 0 0 0 lvtn.3b
flabel comment s 4412 616 4412 616 0 FreeSans 560 0 0 0 lvtn.3a
flabel comment s 3302 -1112 3302 -1112 0 FreeSans 560 0 0 0 lvtn.3b
flabel comment s 4362 -1124 4362 -1124 0 FreeSans 560 0 0 0 lvtn.3a
<< end >>
