magic
tech sky130A
magscale 1 2
timestamp 1607721650
<< metal3 >>
rect 7582 7586 9707 7592
rect 7582 6972 7588 7586
rect 9701 6972 9707 7586
rect 7582 6966 9707 6972
rect 5196 3236 7321 3242
rect 5196 2616 5202 3236
rect 7315 2616 7321 3236
rect 5196 2610 7321 2616
<< via3 >>
rect 7588 6972 9701 7586
rect 5202 2616 7315 3236
<< metal4 >>
rect 7582 7586 9707 7592
rect 7582 6972 7588 7586
rect 9701 6972 9707 7586
rect 7582 6966 9707 6972
rect 5196 3236 7321 3242
rect 5196 2616 5202 3236
rect 7315 2616 7321 3236
rect 5196 2610 7321 2616
<< properties >>
string FIXED_BBOX 0 -406 15000 39593
<< end >>
