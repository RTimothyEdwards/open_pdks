MACRO sky130_fd_io__top_gpio_ovtv2
  CLASS BLOCK ;
  FOREIGN sky130_fd_io__top_gpio_ovtv2 ;
  ORIGIN 0.400 0.735 ;
  SIZE 141.455 BY 201.490 ;
  PIN VSSIO_Q
    PORT
      LAYER met5 ;
        RECT 138.730 58.335 140.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 58.235 140.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    PORT
      LAYER met5 ;
        RECT 138.730 31.985 140.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 31.885 140.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
  END VSWITCH
  PIN VSSIO
    PORT
      LAYER met5 ;
        RECT 138.730 25.935 140.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730 175.785 140.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.365 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 175.785 140.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 25.835 140.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.365 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
  END VSSIO
  PIN VSSD
    PORT
      LAYER met5 ;
        RECT 138.730 41.685 140.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 41.585 140.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
  END VSSD
  PIN VSSA
    PORT
      LAYER met5 ;
        RECT 138.730 36.840 140.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730 47.735 140.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 2.040 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 51.645 140.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 140.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 140.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 36.735 140.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 2.040 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 1.270 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 1.270 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
  END VSSA
  PIN VDDIO_Q
    PORT
      LAYER met5 ;
        RECT 138.730 64.185 140.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 64.085 140.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
  END VDDIO_Q
  PIN VDDIO
    PORT
      LAYER met5 ;
        RECT 138.730 70.035 140.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730 19.885 140.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 19.785 140.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 70.035 140.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
  END VDDIO
  PIN VDDA
    PORT
      LAYER met5 ;
        RECT 139.035 15.035 140.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.035 14.935 140.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
  END VDDA
  PIN VCCHIB
    PORT
      LAYER met5 ;
        RECT 138.730 2.135 140.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 2.035 140.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
  END VCCHIB
  PIN VCCD
    PORT
      LAYER met5 ;
        RECT 138.730 8.985 140.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 8.885 140.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
  END VCCD
  PIN PAD
    PORT
      LAYER met5 ;
        RECT 17.930 117.530 86.325 162.905 ;
    END
  END PAD
  PIN AMUXBUS_A
    PORT
      LAYER met4 ;
        RECT 48.930 53.125 140.000 56.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 38.675 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    PORT
      LAYER met4 ;
        RECT 99.710 48.365 140.000 51.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 85.865 51.345 ;
    END
  END AMUXBUS_B
  PIN DM[0]
    PORT
      LAYER met3 ;
        RECT 129.125 0.000 129.455 20.955 ;
    END
  END DM[0]
  PIN DM[1]
    PORT
      LAYER met3 ;
        RECT 128.275 0.000 128.605 20.180 ;
    END
  END DM[1]
  PIN DM[2]
    PORT
      LAYER met3 ;
        RECT 108.395 0.000 108.725 20.640 ;
    END
  END DM[2]
  PIN INP_DIS
    PORT
      LAYER met3 ;
        RECT 107.545 0.000 107.875 8.060 ;
    END
  END INP_DIS
  PIN VTRIP_SEL
    PORT
      LAYER met3 ;
        RECT 87.665 0.000 87.995 20.980 ;
    END
  END VTRIP_SEL
  PIN IB_MODE_SEL[0]
    PORT
      LAYER met3 ;
        RECT 86.815 0.000 87.145 20.980 ;
    END
  END IB_MODE_SEL[0]
  PIN IB_MODE_SEL[1]
    PORT
      LAYER met3 ;
        RECT 66.935 0.000 67.265 20.980 ;
    END
  END IB_MODE_SEL[1]
  PIN SLEW_CTL[0]
    PORT
      LAYER met3 ;
        RECT 66.085 0.000 66.415 20.980 ;
    END
  END SLEW_CTL[0]
  PIN SLEW_CTL[1]
    PORT
      LAYER met3 ;
        RECT 46.205 0.000 46.535 20.980 ;
    END
  END SLEW_CTL[1]
  PIN HYS_TRIM
    PORT
      LAYER met3 ;
        RECT 45.355 0.000 45.685 8.060 ;
    END
  END HYS_TRIM
  PIN HLD_OVR
    PORT
      LAYER met3 ;
        RECT 27.355 0.000 27.685 14.055 ;
    END
  END HLD_OVR
  PIN ENABLE_H
    PORT
      LAYER met3 ;
        RECT 22.135 0.000 22.465 30.150 ;
    END
  END ENABLE_H
  PIN HLD_H_N
    PORT
      LAYER met3 ;
        RECT 19.635 0.000 19.965 17.985 ;
    END
  END HLD_H_N
  PIN ENABLE_VDDA_H
    PORT
      LAYER met3 ;
        RECT 8.770 0.000 9.100 7.915 ;
    END
  END ENABLE_VDDA_H
  PIN ANALOG_EN
    PORT
      LAYER met3 ;
        RECT 8.115 0.000 8.445 14.070 ;
    END
  END ANALOG_EN
  PIN ENABLE_INP_H
    PORT
      LAYER met3 ;
        RECT 7.110 0.000 7.440 0.670 ;
    END
  END ENABLE_INP_H
  PIN IN
    PORT
      LAYER met3 ;
        RECT 20.380 0.000 20.710 11.310 ;
    END
  END IN
  PIN IN_H
    PORT
      LAYER met3 ;
        RECT 24.380 0.000 24.710 0.940 ;
    END
  END IN_H
  PIN VINREF
    PORT
      LAYER met3 ;
        RECT 44.035 0.000 44.365 4.885 ;
    END
  END VINREF
  PIN OUT
    PORT
      LAYER met3 ;
        RECT 74.125 0.000 74.455 14.865 ;
    END
  END OUT
  PIN ANALOG_POL
    PORT
      LAYER met3 ;
        RECT 65.235 0.000 65.565 1.165 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    PORT
      LAYER met3 ;
        RECT 51.655 0.000 51.985 8.060 ;
    END
  END ANALOG_SEL
  PIN SLOW
    PORT
      LAYER met3 ;
        RECT 125.140 0.000 125.470 11.965 ;
    END
  END SLOW
  PIN OE_N
    PORT
      LAYER met3 ;
        RECT 124.445 0.000 124.775 8.060 ;
    END
  END OE_N
  PIN TIE_HI_ESD
    PORT
      LAYER met3 ;
        RECT 129.975 0.000 130.305 61.655 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    PORT
      LAYER met3 ;
        RECT 115.290 0.000 115.890 39.035 ;
    END
  END TIE_LO_ESD
  PIN PAD_A_ESD_0_H
    PORT
      LAYER met3 ;
        RECT 1.600 0.000 2.200 5.470 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    PORT
      LAYER met3 ;
        RECT 0.330 0.000 0.930 71.380 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    PORT
      LAYER met3 ;
        RECT 2.885 0.000 3.485 5.900 ;
    END
  END PAD_A_NOESD_H
  PIN ENABLE_VSWITCH_H
    PORT
      LAYER met3 ;
        RECT 5.765 0.000 6.365 12.470 ;
    END
  END ENABLE_VSWITCH_H
  PIN ENABLE_VDDIO
    PORT
      LAYER met3 ;
        RECT 95.845 0.000 96.215 20.755 ;
    END
  END ENABLE_VDDIO
  OBS
      LAYER nwell ;
        RECT -0.400 10.495 11.880 11.925 ;
        RECT -0.400 1.430 1.030 10.495 ;
        RECT -0.400 0.000 11.880 1.430 ;
      LAYER li1 ;
        RECT 0.230 0.200 140.475 199.780 ;
      LAYER met1 ;
        RECT 0.080 0.000 140.475 199.810 ;
      LAYER met2 ;
        RECT 0.080 0.000 140.325 199.955 ;
      LAYER met3 ;
        RECT 0.330 71.780 140.000 199.715 ;
        RECT 1.330 62.055 140.000 71.780 ;
        RECT 1.330 39.435 129.575 62.055 ;
        RECT 1.330 30.550 114.890 39.435 ;
        RECT 1.330 18.385 21.735 30.550 ;
        RECT 1.330 14.470 19.235 18.385 ;
        RECT 1.330 12.870 7.715 14.470 ;
        RECT 1.330 6.300 5.365 12.870 ;
        RECT 1.330 5.870 2.485 6.300 ;
        RECT 3.885 0.000 5.365 6.300 ;
        RECT 6.765 1.070 7.715 12.870 ;
        RECT 8.845 8.315 19.235 14.470 ;
        RECT 20.365 11.710 21.735 18.385 ;
        RECT 9.500 0.000 19.235 8.315 ;
        RECT 21.110 0.000 21.735 11.710 ;
        RECT 22.865 21.380 114.890 30.550 ;
        RECT 22.865 14.455 45.805 21.380 ;
        RECT 22.865 1.340 26.955 14.455 ;
        RECT 22.865 0.000 23.980 1.340 ;
        RECT 25.110 0.000 26.955 1.340 ;
        RECT 28.085 8.460 45.805 14.455 ;
        RECT 46.935 8.460 65.685 21.380 ;
        RECT 28.085 5.285 44.955 8.460 ;
        RECT 28.085 0.000 43.635 5.285 ;
        RECT 44.765 0.000 44.955 5.285 ;
        RECT 46.935 0.000 51.255 8.460 ;
        RECT 52.385 1.565 65.685 8.460 ;
        RECT 67.665 15.265 86.415 21.380 ;
        RECT 52.385 0.000 64.835 1.565 ;
        RECT 67.665 0.000 73.725 15.265 ;
        RECT 74.855 0.000 86.415 15.265 ;
        RECT 88.395 21.155 114.890 21.380 ;
        RECT 88.395 0.000 95.445 21.155 ;
        RECT 96.615 21.040 114.890 21.155 ;
        RECT 96.615 8.460 107.995 21.040 ;
        RECT 96.615 0.000 107.145 8.460 ;
        RECT 109.125 0.000 114.890 21.040 ;
        RECT 116.290 21.355 129.575 39.435 ;
        RECT 116.290 20.580 128.725 21.355 ;
        RECT 116.290 12.365 127.875 20.580 ;
        RECT 116.290 8.460 124.740 12.365 ;
        RECT 116.290 0.000 124.045 8.460 ;
        RECT 125.870 0.000 127.875 12.365 ;
        RECT 130.705 0.000 140.000 62.055 ;
      LAYER met4 ;
        RECT 1.765 175.385 138.330 200.000 ;
        RECT 0.965 95.400 139.035 175.385 ;
        RECT 1.670 69.635 138.330 95.400 ;
        RECT 0.965 68.935 139.035 69.635 ;
        RECT 1.670 63.685 138.330 68.935 ;
        RECT 0.965 63.085 139.035 63.685 ;
        RECT 1.670 57.835 138.330 63.085 ;
        RECT 0.965 57.135 139.035 57.835 ;
        RECT 39.075 52.725 48.530 56.005 ;
        RECT 2.440 51.745 138.330 52.725 ;
        RECT 86.265 48.465 99.310 51.745 ;
        RECT 0.965 46.635 139.035 47.335 ;
        RECT 1.670 41.185 138.330 46.635 ;
        RECT 0.965 40.585 139.035 41.185 ;
        RECT 1.670 36.335 138.330 40.585 ;
        RECT 0.965 35.735 139.035 36.335 ;
        RECT 1.670 31.485 138.330 35.735 ;
        RECT 0.965 30.885 139.035 31.485 ;
        RECT 1.670 25.435 138.330 30.885 ;
        RECT 0.965 24.835 139.035 25.435 ;
        RECT 1.670 19.385 138.330 24.835 ;
        RECT 0.965 18.785 139.035 19.385 ;
        RECT 1.365 14.535 138.635 18.785 ;
        RECT 0.965 13.935 139.035 14.535 ;
        RECT 1.670 8.485 138.330 13.935 ;
        RECT 0.965 7.885 139.035 8.485 ;
        RECT 1.670 1.635 138.330 7.885 ;
        RECT 0.965 1.160 139.035 1.635 ;
      LAYER met5 ;
        RECT 2.965 174.185 137.130 200.000 ;
        RECT 0.000 164.505 140.000 174.185 ;
        RECT 0.000 115.930 16.330 164.505 ;
        RECT 87.925 115.930 140.000 164.505 ;
        RECT 0.000 96.585 140.000 115.930 ;
        RECT 2.870 58.335 137.130 96.585 ;
        RECT 3.640 46.135 137.130 58.335 ;
        RECT 2.870 18.285 137.130 46.135 ;
        RECT 2.565 15.035 137.435 18.285 ;
        RECT 2.870 2.135 137.130 15.035 ;
  END
END sky130_fd_io__top_gpio_ovtv2
END LIBRARY

