magic
tech sky130A
magscale 1 2
timestamp 1602972891
<< error_p >>
rect 1419 2270 1664 2276
rect 2097 2235 2343 2239
rect 3033 2229 3045 2235
rect 3055 2229 3067 2235
rect 2096 2207 2342 2211
rect 2679 2183 2681 2217
rect 2711 2183 2713 2217
rect 3021 2211 3027 2223
rect 3073 2211 3079 2223
rect 3554 2208 3588 2242
rect 3995 2214 4032 2254
rect 1407 1398 1449 1423
rect 1407 1342 1449 1367
rect 3303 1040 3320 1367
<< locali >>
rect 2665 2217 2733 2239
rect 2665 2183 2679 2217
rect 2713 2183 2733 2217
rect 2665 2172 2733 2183
rect 3019 2223 3087 2245
rect 3019 2189 3033 2223
rect 3067 2189 3087 2223
rect 3019 2178 3087 2189
<< viali >>
rect 2679 2183 2713 2217
rect 3033 2189 3067 2223
<< metal1 >>
rect 1419 2248 1664 2270
rect 2097 2235 2343 2272
rect 2675 2217 2717 2258
rect 3950 2254 4077 2299
rect 2096 2174 2342 2211
rect 2675 2183 2679 2217
rect 2713 2183 2717 2217
rect 2675 2160 2717 2183
rect 3027 2223 3073 2229
rect 3027 2189 3033 2223
rect 3067 2189 3073 2223
rect 3554 2208 3588 2242
rect 3950 2214 3995 2254
rect 4032 2214 4077 2254
rect 3027 2148 3073 2189
rect 3950 2169 4077 2214
rect 1449 1433 2149 1583
rect 1407 1398 2149 1433
rect 1449 1367 2149 1398
rect 1407 1332 2149 1367
rect 1449 883 2149 1332
rect 2564 866 3264 1566
rect 3303 1040 3332 1367
<< labels >>
flabel comment s 500 1677 500 1677 0 FreeSans 560 0 0 0 Not implemented
flabel comment s 1549 2081 1549 2081 0 FreeSans 560 0 0 0 m1.1
flabel comment s 2260 2050 2260 2050 0 FreeSans 560 0 0 0 m1.2
flabel comment s 1821 811 1821 811 0 FreeSans 560 0 0 0 m1.3a
flabel comment s 2974 811 2974 811 0 FreeSans 560 0 0 0 m1.3b
flabel comment s 2708 2080 2708 2080 0 FreeSans 560 0 0 0 m1.4
flabel comment s 568 1459 568 1459 0 FreeSans 560 0 0 0 m1.4a
flabel comment s 3061 2094 3061 2094 0 FreeSans 560 0 0 0 m1.5
flabel comment s 3599 2100 3599 2100 0 FreeSans 560 0 0 0 m1.6
flabel comment s 3991 2098 3991 2098 0 FreeSans 560 0 0 0 m1.7
flabel comment s 493 2348 493 2348 0 FreeSans 800 0 0 0 Met1 (m1)
<< end >>
