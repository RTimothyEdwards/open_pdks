magic
tech sky130A
magscale 1 2
timestamp 1602597384
<< error_s >>
rect 308 39412 2226 39494
rect 95 38277 177 39311
rect 387 38447 469 39141
rect 609 39130 1915 39212
rect 777 38936 1719 38986
rect 646 38893 672 38904
rect 662 38853 756 38893
rect 1668 38853 1762 38893
rect 662 38693 756 38733
rect 1668 38693 1762 38733
rect 646 38682 672 38693
rect 777 38592 1719 38642
rect 609 38378 1915 38460
rect 1955 38447 2037 39141
rect 2247 38277 2329 39311
rect 3148 38410 3198 39410
rect 3298 38410 3426 39410
rect 3454 38410 3504 39410
rect 3570 38410 3620 39410
rect 3780 38410 3836 39410
rect 3996 38410 4052 39410
rect 4152 38410 4280 39410
rect 4308 38410 4358 39410
rect 4474 38410 4524 39410
rect 4684 38410 4740 39410
rect 4840 38410 4968 39410
rect 4996 38410 5052 39410
rect 5152 38410 5280 39410
rect 5308 38410 5364 39410
rect 5464 38410 5514 39410
rect 5580 38410 5630 39010
rect 5730 38410 5780 39010
rect 5846 38410 5896 39410
rect 5996 38410 6052 39410
rect 6152 38410 6202 39410
rect 7092 38406 7150 38440
rect 7932 38418 7982 39418
rect 8082 38418 8210 39418
rect 8238 38418 8366 39418
rect 8394 38418 8522 39418
rect 8550 38418 8678 39418
rect 8706 38418 8756 39418
rect 8822 38418 8872 39418
rect 8972 38418 9028 39418
rect 9128 38418 9178 39418
rect 9244 38418 9294 39418
rect 9394 38418 9522 39418
rect 9550 38418 9606 39418
rect 9706 38418 9834 39418
rect 9862 38418 9912 39418
rect 9978 38418 10028 39418
rect 10128 38418 10256 39418
rect 10284 38418 10340 39418
rect 10440 38418 10568 39418
rect 10596 38790 10646 39418
rect 10596 38718 10649 38790
rect 10596 38418 10646 38718
rect 10709 38418 10721 38718
rect 14297 38255 15297 38305
rect 2355 38203 2358 38204
rect 2355 38202 2356 38203
rect 2357 38202 2358 38203
rect 2355 38201 2358 38202
rect 308 38093 2226 38175
rect 14297 38099 15297 38227
rect 2355 38066 2358 38067
rect 2355 38065 2356 38066
rect 2357 38065 2358 38066
rect 2355 38064 2358 38065
rect 95 36957 177 37991
rect 387 37127 469 37821
rect 609 37808 1915 37890
rect 777 37626 1719 37676
rect 646 37575 672 37586
rect 662 37553 756 37575
rect 662 37535 672 37553
rect 694 37535 756 37553
rect 1668 37553 1762 37575
rect 1668 37535 1730 37553
rect 1752 37535 1762 37553
rect 662 37397 672 37415
rect 694 37397 756 37415
rect 662 37375 756 37397
rect 1668 37397 1730 37415
rect 1752 37397 1762 37415
rect 1668 37375 1762 37397
rect 646 37364 672 37375
rect 777 37282 1719 37332
rect 609 37056 1915 37138
rect 1955 37127 2037 37821
rect 2247 36957 2329 37991
rect 8191 37965 9191 38015
rect 9587 37965 10187 38015
rect 8191 37809 9191 37937
rect 11931 37905 12931 37955
rect 14297 37949 15297 37999
rect 9587 37809 10187 37865
rect 8191 37653 9191 37781
rect 9587 37653 10187 37709
rect 11931 37689 12931 37817
rect 8191 37503 9191 37553
rect 9587 37497 10187 37553
rect 11931 37479 12931 37529
rect 9587 37347 10187 37397
rect 308 36774 2226 36856
rect 1021 36719 1191 36774
rect 2255 36719 2424 36787
rect 1089 36679 1191 36719
rect 2323 36679 2424 36719
rect 1089 36638 1123 36679
rect 2323 36638 2357 36679
rect 1398 36418 1998 36468
rect 1398 36168 1998 36218
rect 3118 35743 3168 36743
rect 3328 35743 3456 36743
rect 3544 35743 3672 36743
rect 3760 35743 3888 36743
rect 3976 35743 4104 36743
rect 4192 35743 4248 36743
rect 4408 35743 4464 36743
rect 4624 35743 4752 36743
rect 4840 35743 4968 36743
rect 5056 35743 5184 36743
rect 5272 35743 5400 36743
rect 5488 35743 5544 36743
rect 5704 35743 5832 36743
rect 5920 35743 6048 36743
rect 6136 35743 6264 36743
rect 6352 35743 6402 36743
rect 6468 35743 6518 36743
rect 6678 35743 6728 36743
rect 6794 35743 6844 36743
rect 7004 35743 7054 36743
rect 7120 35743 7170 36743
rect 7330 35743 7380 36743
rect 7443 36558 7455 36758
rect 7446 35743 7496 36343
rect 7696 35743 7752 36343
rect 7852 35743 7980 36343
rect 8008 35743 8064 36343
rect 8164 35743 8292 36343
rect 8320 35743 8370 36343
rect 8436 35743 8486 36743
rect 8586 35743 8642 36743
rect 8742 35743 8792 36743
rect 8870 35743 8920 36743
rect 9020 35743 9148 36743
rect 9176 35743 9304 36743
rect 9332 35743 9388 36743
rect 9488 35743 9616 36743
rect 9644 35743 9772 36743
rect 9800 35743 9928 36743
rect 9956 35743 10006 36743
rect 10072 35743 10122 36743
rect 10222 35743 10350 36743
rect 10378 35743 10506 36743
rect 10534 35743 10662 36743
rect 10690 35743 10746 36743
rect 10846 35743 10974 36743
rect 11002 35743 11130 36743
rect 11158 35743 11214 36743
rect 11314 35743 11364 36743
rect 12585 36543 12638 36743
rect 12588 35743 12638 36543
rect 12798 35743 12926 36743
rect 13014 35743 13070 36743
rect 13230 35743 13358 36743
rect 13446 35743 13496 36743
rect 13562 35743 13612 36743
rect 13772 35743 13822 36743
rect 11309 35656 11345 35667
rect 11461 35656 13785 35667
rect 11309 35634 13785 35656
rect 11309 35633 11345 35634
rect 11461 35633 13785 35634
rect 6371 34402 13485 34424
rect 1697 34055 2697 34105
rect 2807 34055 3807 34105
rect 3928 34055 4928 34105
rect 5049 34055 6049 34105
rect 6606 34055 7606 34105
rect 7727 34055 8727 34105
rect 8848 34055 9848 34105
rect 9958 34055 10958 34105
rect 11079 34055 12079 34105
rect 12200 34055 13200 34105
rect 1697 33885 2697 33935
rect 2807 33885 3807 33935
rect 3928 33885 4928 33935
rect 5049 33885 6049 33935
rect 6606 33885 7606 33935
rect 7727 33885 8727 33935
rect 8848 33885 9848 33935
rect 9958 33885 10958 33935
rect 11079 33885 12079 33935
rect 12200 33885 13200 33935
rect 1302 33622 1437 33626
rect 6311 33622 6345 33626
rect 13414 33622 13553 33656
rect 1302 33598 13553 33622
rect 15317 33612 15331 34456
rect 15307 33598 15331 33612
rect 1302 33588 15331 33598
rect 1301 33572 15331 33588
rect 1302 33534 13482 33572
rect 13485 33534 13495 33572
rect 1924 32204 2134 32240
rect 14186 32204 14299 32240
rect 14748 32204 15030 32240
rect 1513 31204 1591 32204
rect 1713 31204 1785 32204
rect 1936 31204 1960 32204
rect 2001 31204 2057 32204
rect 2098 31204 2134 32204
rect 2359 31204 2419 32204
rect 2619 31204 2691 32204
rect 2921 31204 2977 32204
rect 2993 31204 3049 32204
rect 3351 31204 3411 32204
rect 3611 31204 3683 32204
rect 3913 31204 3969 32204
rect 3985 31204 4041 32204
rect 4343 31204 4403 32204
rect 4603 31204 4675 32204
rect 4905 31204 4961 32204
rect 4977 31204 5033 32204
rect 5335 31204 5395 32204
rect 5595 31204 5667 32204
rect 5897 31204 5953 32204
rect 5969 31204 6025 32204
rect 6327 31204 6387 32204
rect 6587 31204 6659 32204
rect 6889 31204 6945 32204
rect 6961 31204 7017 32204
rect 7319 31204 7379 32204
rect 7579 31204 7651 32204
rect 7881 31204 7937 32204
rect 7953 31204 8009 32204
rect 8311 31204 8371 32204
rect 8571 31204 8643 32204
rect 8873 31204 8929 32204
rect 8945 31204 9001 32204
rect 9303 31204 9363 32204
rect 9563 31204 9635 32204
rect 9865 31204 9921 32204
rect 9937 31204 9993 32204
rect 10295 31204 10355 32204
rect 10555 31204 10627 32204
rect 10857 31204 10913 32204
rect 10929 31204 10985 32204
rect 11287 31204 11347 32204
rect 11547 31204 11619 32204
rect 11849 31204 11905 32204
rect 11921 31204 11977 32204
rect 12279 31204 12339 32204
rect 12539 31204 12611 32204
rect 12841 31204 12897 32204
rect 12913 31204 12969 32204
rect 13271 31204 13331 32204
rect 13531 31204 13603 32204
rect 13833 31204 13889 32204
rect 13905 31204 13961 32204
rect 14186 31204 14222 32204
rect 14263 31204 14299 32204
rect 14523 31204 14595 32204
rect 14748 31204 14784 32204
rect 14825 31204 14881 32204
rect 14897 31204 14953 32204
rect 14994 31204 15030 32204
rect 15241 31204 15301 32204
rect 15337 32187 15441 32204
rect 15337 32153 15431 32187
rect 15441 32153 15475 32187
rect 15337 32116 15441 32153
rect 15337 32082 15431 32116
rect 15441 32082 15475 32116
rect 15337 32042 15441 32082
rect 15337 32008 15431 32042
rect 15441 32008 15475 32042
rect 15337 31971 15441 32008
rect 15337 31937 15431 31971
rect 15441 31937 15475 31971
rect 15337 31897 15441 31937
rect 15337 31863 15431 31897
rect 15441 31863 15475 31897
rect 15337 31826 15441 31863
rect 15337 31792 15431 31826
rect 15441 31792 15475 31826
rect 15337 31752 15441 31792
rect 15337 31718 15431 31752
rect 15441 31718 15475 31752
rect 15337 31681 15441 31718
rect 15337 31647 15431 31681
rect 15441 31647 15475 31681
rect 15337 31607 15441 31647
rect 15337 31573 15431 31607
rect 15441 31573 15475 31607
rect 15337 31536 15441 31573
rect 15337 31502 15431 31536
rect 15441 31502 15475 31536
rect 15337 31462 15441 31502
rect 15337 31428 15431 31462
rect 15441 31428 15475 31462
rect 15337 31391 15441 31428
rect 15337 31357 15431 31391
rect 15441 31357 15475 31391
rect 15337 31297 15441 31357
rect 15337 31263 15431 31297
rect 15441 31263 15475 31297
rect 15337 31227 15441 31263
rect 15337 31204 15465 31227
rect 1924 31168 2134 31204
rect 14186 31168 14299 31204
rect 14748 31168 15030 31204
rect 1479 30631 1523 30637
rect 1479 30603 1489 30631
rect 1513 30603 1523 30631
rect 1924 30603 2134 30639
rect 14186 30603 14299 30639
rect 14748 30603 15030 30639
rect 15431 30603 15441 30627
rect 1513 29603 1617 30603
rect 1713 29603 1785 30603
rect 1959 29603 1960 30603
rect 2001 29603 2057 30603
rect 2098 29603 2099 30603
rect 2359 29603 2419 30603
rect 2619 29603 2691 30603
rect 2921 29603 2977 30603
rect 2993 29603 3049 30603
rect 3351 29603 3411 30603
rect 3611 29603 3683 30603
rect 3913 29603 3969 30603
rect 3985 29603 4041 30603
rect 4343 29603 4403 30603
rect 4603 29603 4675 30603
rect 4905 29603 4961 30603
rect 4977 29603 5033 30603
rect 5335 29603 5395 30603
rect 5595 29603 5667 30603
rect 5897 29603 5953 30603
rect 5969 29603 6025 30603
rect 6327 29603 6387 30603
rect 6587 29603 6659 30603
rect 6889 29603 6945 30603
rect 6961 29603 7017 30603
rect 7319 29603 7379 30603
rect 7579 29603 7651 30603
rect 7881 29603 7937 30603
rect 7953 29603 8009 30603
rect 8311 29603 8371 30603
rect 8571 29603 8643 30603
rect 8873 29603 8929 30603
rect 8945 29603 9001 30603
rect 9303 29603 9363 30603
rect 9563 29603 9635 30603
rect 9865 29603 9921 30603
rect 9937 29603 9993 30603
rect 10295 29603 10355 30603
rect 10555 29603 10627 30603
rect 10857 29603 10913 30603
rect 10929 29603 10985 30603
rect 11287 29603 11347 30603
rect 11547 29603 11619 30603
rect 11849 29603 11905 30603
rect 11921 29603 11977 30603
rect 12279 29603 12339 30603
rect 12539 29603 12611 30603
rect 12841 29603 12897 30603
rect 12913 29603 12969 30603
rect 13271 29603 13331 30603
rect 13531 29603 13603 30603
rect 13833 29603 13889 30603
rect 13905 29603 13961 30603
rect 14186 29603 14222 30603
rect 14263 29603 14299 30603
rect 14523 29603 14595 30603
rect 14748 29603 14784 30603
rect 14825 29603 14881 30603
rect 14897 29603 14953 30603
rect 14994 29603 15030 30603
rect 15241 29603 15301 30603
rect 15337 30581 15431 30603
rect 15441 30581 15465 30603
rect 15337 30547 15441 30581
rect 15337 30513 15431 30547
rect 15441 30513 15465 30547
rect 15337 30473 15441 30513
rect 15337 30439 15431 30473
rect 15441 30439 15475 30473
rect 15337 30396 15441 30439
rect 15337 30362 15431 30396
rect 15441 30362 15475 30396
rect 15337 30302 15441 30362
rect 15337 30268 15431 30302
rect 15441 30268 15475 30302
rect 15337 30231 15441 30268
rect 15337 30197 15431 30231
rect 15441 30197 15475 30231
rect 15337 30157 15441 30197
rect 15337 30123 15431 30157
rect 15441 30123 15475 30157
rect 15337 30086 15441 30123
rect 15337 30052 15431 30086
rect 15441 30052 15475 30086
rect 15337 30012 15441 30052
rect 15337 29978 15431 30012
rect 15441 29978 15475 30012
rect 15337 29941 15441 29978
rect 15337 29907 15431 29941
rect 15441 29907 15475 29941
rect 15337 29867 15441 29907
rect 15337 29833 15431 29867
rect 15441 29833 15475 29867
rect 15337 29796 15441 29833
rect 15337 29762 15431 29796
rect 15441 29762 15475 29796
rect 15337 29722 15441 29762
rect 15337 29688 15431 29722
rect 15441 29688 15475 29722
rect 15337 29651 15441 29688
rect 15337 29617 15431 29651
rect 15441 29617 15475 29651
rect 15337 29603 15441 29617
rect 1924 29567 2134 29603
rect 14186 29567 14299 29603
rect 14748 29567 15030 29603
rect 1336 27100 1352 27166
rect 3360 27100 3376 27166
rect 9527 27034 9543 27050
rect 9425 26728 9543 27034
rect 9527 26712 9543 26728
rect 11715 27034 11731 27050
rect 11715 26728 11833 27034
rect 11715 26712 11731 26728
rect 959 24846 983 25638
rect 828 24749 983 24846
rect 828 20203 935 24749
rect 1623 22915 1673 23915
rect 1884 22915 1940 23915
rect 1956 22915 2012 23915
rect 2314 23835 2514 23915
rect 2529 23845 2563 23869
rect 2574 23845 2646 23915
rect 2529 23835 2646 23845
rect 2301 23811 2646 23835
rect 2314 23767 2514 23811
rect 2529 23801 2553 23811
rect 2529 23777 2563 23801
rect 2574 23777 2646 23811
rect 2529 23767 2646 23777
rect 2301 23743 2646 23767
rect 2314 23699 2514 23743
rect 2529 23733 2553 23743
rect 2529 23709 2563 23733
rect 2574 23709 2646 23743
rect 2529 23699 2646 23709
rect 2301 23675 2646 23699
rect 2314 23631 2514 23675
rect 2529 23665 2553 23675
rect 2529 23641 2563 23665
rect 2574 23641 2646 23675
rect 2529 23631 2646 23641
rect 2301 23607 2646 23631
rect 2314 23563 2514 23607
rect 2529 23597 2553 23607
rect 2529 23573 2563 23597
rect 2574 23573 2646 23607
rect 2529 23563 2646 23573
rect 2301 23539 2646 23563
rect 2314 23495 2514 23539
rect 2529 23529 2553 23539
rect 2529 23505 2563 23529
rect 2574 23505 2646 23539
rect 2529 23495 2646 23505
rect 2301 23471 2646 23495
rect 2314 23427 2514 23471
rect 2529 23461 2553 23471
rect 2529 23437 2563 23461
rect 2574 23437 2646 23471
rect 2529 23427 2646 23437
rect 2301 23403 2646 23427
rect 2314 23359 2514 23403
rect 2529 23393 2553 23403
rect 2529 23369 2563 23393
rect 2574 23369 2646 23403
rect 2529 23359 2646 23369
rect 2301 23335 2646 23359
rect 2314 23291 2514 23335
rect 2529 23325 2553 23335
rect 2529 23301 2563 23325
rect 2574 23301 2646 23335
rect 2529 23291 2646 23301
rect 2301 23267 2646 23291
rect 2314 23223 2514 23267
rect 2529 23257 2553 23267
rect 2529 23233 2563 23257
rect 2574 23233 2646 23267
rect 2529 23223 2646 23233
rect 2301 23199 2646 23223
rect 2314 23155 2514 23199
rect 2529 23189 2553 23199
rect 2529 23165 2563 23189
rect 2574 23165 2646 23199
rect 2529 23155 2646 23165
rect 2301 23131 2646 23155
rect 2314 23087 2514 23131
rect 2529 23121 2553 23131
rect 2529 23097 2563 23121
rect 2574 23097 2646 23131
rect 2529 23087 2646 23097
rect 2301 23063 2646 23087
rect 2314 23019 2514 23063
rect 2529 23053 2553 23063
rect 2529 23029 2563 23053
rect 2574 23029 2646 23063
rect 2529 23019 2646 23029
rect 2301 22995 2646 23019
rect 2314 22951 2514 22995
rect 2529 22985 2553 22995
rect 2529 22961 2563 22985
rect 2574 22961 2646 22995
rect 2529 22951 2646 22961
rect 2301 22927 2646 22951
rect 2314 22915 2514 22927
rect 2325 22903 2349 22915
rect 2529 22903 2553 22927
rect 2574 22915 2646 22927
rect 2876 22915 2932 23915
rect 2948 22915 3004 23915
rect 3306 23835 3506 23915
rect 3521 23845 3555 23869
rect 3566 23845 3638 23915
rect 3521 23835 3638 23845
rect 3293 23811 3638 23835
rect 3306 23767 3506 23811
rect 3521 23801 3545 23811
rect 3521 23777 3555 23801
rect 3566 23777 3638 23811
rect 3521 23767 3638 23777
rect 3293 23743 3638 23767
rect 3306 23699 3506 23743
rect 3521 23733 3545 23743
rect 3521 23709 3555 23733
rect 3566 23709 3638 23743
rect 3521 23699 3638 23709
rect 3293 23675 3638 23699
rect 3306 23631 3506 23675
rect 3521 23665 3545 23675
rect 3521 23641 3555 23665
rect 3566 23641 3638 23675
rect 3521 23631 3638 23641
rect 3293 23607 3638 23631
rect 3306 23563 3506 23607
rect 3521 23597 3545 23607
rect 3521 23573 3555 23597
rect 3566 23573 3638 23607
rect 3521 23563 3638 23573
rect 3293 23539 3638 23563
rect 3306 23495 3506 23539
rect 3521 23529 3545 23539
rect 3521 23505 3555 23529
rect 3566 23505 3638 23539
rect 3521 23495 3638 23505
rect 3293 23471 3638 23495
rect 3306 23427 3506 23471
rect 3521 23461 3545 23471
rect 3521 23437 3555 23461
rect 3566 23437 3638 23471
rect 3521 23427 3638 23437
rect 3293 23403 3638 23427
rect 3306 23359 3506 23403
rect 3521 23393 3545 23403
rect 3521 23369 3555 23393
rect 3566 23369 3638 23403
rect 3521 23359 3638 23369
rect 3293 23335 3638 23359
rect 3306 23291 3506 23335
rect 3521 23325 3545 23335
rect 3521 23301 3555 23325
rect 3566 23301 3638 23335
rect 3521 23291 3638 23301
rect 3293 23267 3638 23291
rect 3306 23223 3506 23267
rect 3521 23257 3545 23267
rect 3521 23233 3555 23257
rect 3566 23233 3638 23267
rect 3521 23223 3638 23233
rect 3293 23199 3638 23223
rect 3306 23155 3506 23199
rect 3521 23189 3545 23199
rect 3521 23165 3555 23189
rect 3566 23165 3638 23199
rect 3521 23155 3638 23165
rect 3293 23131 3638 23155
rect 3306 23087 3506 23131
rect 3521 23121 3545 23131
rect 3521 23097 3555 23121
rect 3566 23097 3638 23131
rect 3521 23087 3638 23097
rect 3293 23063 3638 23087
rect 3306 23019 3506 23063
rect 3521 23053 3545 23063
rect 3521 23029 3555 23053
rect 3566 23029 3638 23063
rect 3521 23019 3638 23029
rect 3293 22995 3638 23019
rect 3306 22951 3506 22995
rect 3521 22985 3545 22995
rect 3521 22961 3555 22985
rect 3566 22961 3638 22995
rect 3521 22951 3638 22961
rect 3293 22927 3638 22951
rect 3306 22915 3506 22927
rect 3317 22903 3341 22915
rect 3521 22903 3545 22927
rect 3566 22915 3638 22927
rect 3868 22915 3924 23915
rect 3940 22915 3996 23915
rect 4298 23835 4498 23915
rect 4513 23845 4547 23869
rect 4558 23845 4630 23915
rect 4513 23835 4630 23845
rect 4285 23811 4630 23835
rect 4298 23767 4498 23811
rect 4513 23801 4537 23811
rect 4513 23777 4547 23801
rect 4558 23777 4630 23811
rect 4513 23767 4630 23777
rect 4285 23743 4630 23767
rect 4298 23699 4498 23743
rect 4513 23733 4537 23743
rect 4513 23709 4547 23733
rect 4558 23709 4630 23743
rect 4513 23699 4630 23709
rect 4285 23675 4630 23699
rect 4298 23631 4498 23675
rect 4513 23665 4537 23675
rect 4513 23641 4547 23665
rect 4558 23641 4630 23675
rect 4513 23631 4630 23641
rect 4285 23607 4630 23631
rect 4298 23563 4498 23607
rect 4513 23597 4537 23607
rect 4513 23573 4547 23597
rect 4558 23573 4630 23607
rect 4513 23563 4630 23573
rect 4285 23539 4630 23563
rect 4298 23495 4498 23539
rect 4513 23529 4537 23539
rect 4513 23505 4547 23529
rect 4558 23505 4630 23539
rect 4513 23495 4630 23505
rect 4285 23471 4630 23495
rect 4298 23427 4498 23471
rect 4513 23461 4537 23471
rect 4513 23437 4547 23461
rect 4558 23437 4630 23471
rect 4513 23427 4630 23437
rect 4285 23403 4630 23427
rect 4298 23359 4498 23403
rect 4513 23393 4537 23403
rect 4513 23369 4547 23393
rect 4558 23369 4630 23403
rect 4513 23359 4630 23369
rect 4285 23335 4630 23359
rect 4298 23291 4498 23335
rect 4513 23325 4537 23335
rect 4513 23301 4547 23325
rect 4558 23301 4630 23335
rect 4513 23291 4630 23301
rect 4285 23267 4630 23291
rect 4298 23223 4498 23267
rect 4513 23257 4537 23267
rect 4513 23233 4547 23257
rect 4558 23233 4630 23267
rect 4513 23223 4630 23233
rect 4285 23199 4630 23223
rect 4298 23155 4498 23199
rect 4513 23189 4537 23199
rect 4513 23165 4547 23189
rect 4558 23165 4630 23199
rect 4513 23155 4630 23165
rect 4285 23131 4630 23155
rect 4298 23087 4498 23131
rect 4513 23121 4537 23131
rect 4513 23097 4547 23121
rect 4558 23097 4630 23131
rect 4513 23087 4630 23097
rect 4285 23063 4630 23087
rect 4298 23019 4498 23063
rect 4513 23053 4537 23063
rect 4513 23029 4547 23053
rect 4558 23029 4630 23063
rect 4513 23019 4630 23029
rect 4285 22995 4630 23019
rect 4298 22951 4498 22995
rect 4513 22985 4537 22995
rect 4513 22961 4547 22985
rect 4558 22961 4630 22995
rect 4513 22951 4630 22961
rect 4285 22927 4630 22951
rect 4298 22915 4498 22927
rect 4309 22903 4333 22915
rect 4513 22903 4537 22927
rect 4558 22915 4630 22927
rect 4860 22915 4916 23915
rect 4932 22915 4988 23915
rect 5290 23835 5490 23915
rect 5505 23845 5539 23869
rect 5550 23845 5622 23915
rect 5505 23835 5622 23845
rect 5277 23811 5622 23835
rect 5290 23767 5490 23811
rect 5505 23801 5529 23811
rect 5505 23777 5539 23801
rect 5550 23777 5622 23811
rect 5505 23767 5622 23777
rect 5277 23743 5622 23767
rect 5290 23699 5490 23743
rect 5505 23733 5529 23743
rect 5505 23709 5539 23733
rect 5550 23709 5622 23743
rect 5505 23699 5622 23709
rect 5277 23675 5622 23699
rect 5290 23631 5490 23675
rect 5505 23665 5529 23675
rect 5505 23641 5539 23665
rect 5550 23641 5622 23675
rect 5505 23631 5622 23641
rect 5277 23607 5622 23631
rect 5290 23563 5490 23607
rect 5505 23597 5529 23607
rect 5505 23573 5539 23597
rect 5550 23573 5622 23607
rect 5505 23563 5622 23573
rect 5277 23539 5622 23563
rect 5290 23495 5490 23539
rect 5505 23529 5529 23539
rect 5505 23505 5539 23529
rect 5550 23505 5622 23539
rect 5505 23495 5622 23505
rect 5277 23471 5622 23495
rect 5290 23427 5490 23471
rect 5505 23461 5529 23471
rect 5505 23437 5539 23461
rect 5550 23437 5622 23471
rect 5505 23427 5622 23437
rect 5277 23403 5622 23427
rect 5290 23359 5490 23403
rect 5505 23393 5529 23403
rect 5505 23369 5539 23393
rect 5550 23369 5622 23403
rect 5505 23359 5622 23369
rect 5277 23335 5622 23359
rect 5290 23291 5490 23335
rect 5505 23325 5529 23335
rect 5505 23301 5539 23325
rect 5550 23301 5622 23335
rect 5505 23291 5622 23301
rect 5277 23267 5622 23291
rect 5290 23223 5490 23267
rect 5505 23257 5529 23267
rect 5505 23233 5539 23257
rect 5550 23233 5622 23267
rect 5505 23223 5622 23233
rect 5277 23199 5622 23223
rect 5290 23155 5490 23199
rect 5505 23189 5529 23199
rect 5505 23165 5539 23189
rect 5550 23165 5622 23199
rect 5505 23155 5622 23165
rect 5277 23131 5622 23155
rect 5290 23087 5490 23131
rect 5505 23121 5529 23131
rect 5505 23097 5539 23121
rect 5550 23097 5622 23131
rect 5505 23087 5622 23097
rect 5277 23063 5622 23087
rect 5290 23019 5490 23063
rect 5505 23053 5529 23063
rect 5505 23029 5539 23053
rect 5550 23029 5622 23063
rect 5505 23019 5622 23029
rect 5277 22995 5622 23019
rect 5290 22951 5490 22995
rect 5505 22985 5529 22995
rect 5505 22961 5539 22985
rect 5550 22961 5622 22995
rect 5505 22951 5622 22961
rect 5277 22927 5622 22951
rect 5290 22915 5490 22927
rect 5301 22903 5325 22915
rect 5505 22903 5529 22927
rect 5550 22915 5622 22927
rect 5852 22915 5908 23915
rect 5924 22915 5980 23915
rect 6282 23835 6482 23915
rect 6497 23845 6531 23869
rect 6542 23845 6614 23915
rect 6497 23835 6614 23845
rect 6269 23811 6614 23835
rect 6282 23767 6482 23811
rect 6497 23801 6521 23811
rect 6497 23777 6531 23801
rect 6542 23777 6614 23811
rect 6497 23767 6614 23777
rect 6269 23743 6614 23767
rect 6282 23699 6482 23743
rect 6497 23733 6521 23743
rect 6497 23709 6531 23733
rect 6542 23709 6614 23743
rect 6497 23699 6614 23709
rect 6269 23675 6614 23699
rect 6282 23631 6482 23675
rect 6497 23665 6521 23675
rect 6497 23641 6531 23665
rect 6542 23641 6614 23675
rect 6497 23631 6614 23641
rect 6269 23607 6614 23631
rect 6282 23563 6482 23607
rect 6497 23597 6521 23607
rect 6497 23573 6531 23597
rect 6542 23573 6614 23607
rect 6497 23563 6614 23573
rect 6269 23539 6614 23563
rect 6282 23495 6482 23539
rect 6497 23529 6521 23539
rect 6497 23505 6531 23529
rect 6542 23505 6614 23539
rect 6497 23495 6614 23505
rect 6269 23471 6614 23495
rect 6282 23427 6482 23471
rect 6497 23461 6521 23471
rect 6497 23437 6531 23461
rect 6542 23437 6614 23471
rect 6497 23427 6614 23437
rect 6269 23403 6614 23427
rect 6282 23359 6482 23403
rect 6497 23393 6521 23403
rect 6497 23369 6531 23393
rect 6542 23369 6614 23403
rect 6497 23359 6614 23369
rect 6269 23335 6614 23359
rect 6282 23291 6482 23335
rect 6497 23325 6521 23335
rect 6497 23301 6531 23325
rect 6542 23301 6614 23335
rect 6497 23291 6614 23301
rect 6269 23267 6614 23291
rect 6282 23223 6482 23267
rect 6497 23257 6521 23267
rect 6497 23233 6531 23257
rect 6542 23233 6614 23267
rect 6497 23223 6614 23233
rect 6269 23199 6614 23223
rect 6282 23155 6482 23199
rect 6497 23189 6521 23199
rect 6497 23165 6531 23189
rect 6542 23165 6614 23199
rect 6497 23155 6614 23165
rect 6269 23131 6614 23155
rect 6282 23087 6482 23131
rect 6497 23121 6521 23131
rect 6497 23097 6531 23121
rect 6542 23097 6614 23131
rect 6497 23087 6614 23097
rect 6269 23063 6614 23087
rect 6282 23019 6482 23063
rect 6497 23053 6521 23063
rect 6497 23029 6531 23053
rect 6542 23029 6614 23063
rect 6497 23019 6614 23029
rect 6269 22995 6614 23019
rect 6282 22951 6482 22995
rect 6497 22985 6521 22995
rect 6497 22961 6531 22985
rect 6542 22961 6614 22995
rect 6497 22951 6614 22961
rect 6269 22927 6614 22951
rect 6282 22915 6482 22927
rect 6293 22903 6317 22915
rect 6497 22903 6521 22927
rect 6542 22915 6614 22927
rect 6844 22915 6900 23915
rect 6916 22915 6972 23915
rect 7274 23835 7474 23915
rect 7489 23845 7523 23869
rect 7534 23845 7606 23915
rect 7489 23835 7606 23845
rect 7261 23811 7606 23835
rect 7274 23767 7474 23811
rect 7489 23801 7513 23811
rect 7489 23777 7523 23801
rect 7534 23777 7606 23811
rect 7489 23767 7606 23777
rect 7261 23743 7606 23767
rect 7274 23699 7474 23743
rect 7489 23733 7513 23743
rect 7489 23709 7523 23733
rect 7534 23709 7606 23743
rect 7489 23699 7606 23709
rect 7261 23675 7606 23699
rect 7274 23631 7474 23675
rect 7489 23665 7513 23675
rect 7489 23641 7523 23665
rect 7534 23641 7606 23675
rect 7489 23631 7606 23641
rect 7261 23607 7606 23631
rect 7274 23563 7474 23607
rect 7489 23597 7513 23607
rect 7489 23573 7523 23597
rect 7534 23573 7606 23607
rect 7489 23563 7606 23573
rect 7261 23539 7606 23563
rect 7274 23495 7474 23539
rect 7489 23529 7513 23539
rect 7489 23505 7523 23529
rect 7534 23505 7606 23539
rect 7489 23495 7606 23505
rect 7261 23471 7606 23495
rect 7274 23427 7474 23471
rect 7489 23461 7513 23471
rect 7489 23437 7523 23461
rect 7534 23437 7606 23471
rect 7489 23427 7606 23437
rect 7261 23403 7606 23427
rect 7274 23359 7474 23403
rect 7489 23393 7513 23403
rect 7489 23369 7523 23393
rect 7534 23369 7606 23403
rect 7489 23359 7606 23369
rect 7261 23335 7606 23359
rect 7274 23291 7474 23335
rect 7489 23325 7513 23335
rect 7489 23301 7523 23325
rect 7534 23301 7606 23335
rect 7489 23291 7606 23301
rect 7261 23267 7606 23291
rect 7274 23223 7474 23267
rect 7489 23257 7513 23267
rect 7489 23233 7523 23257
rect 7534 23233 7606 23267
rect 7489 23223 7606 23233
rect 7261 23199 7606 23223
rect 7274 23155 7474 23199
rect 7489 23189 7513 23199
rect 7489 23165 7523 23189
rect 7534 23165 7606 23199
rect 7489 23155 7606 23165
rect 7261 23131 7606 23155
rect 7274 23087 7474 23131
rect 7489 23121 7513 23131
rect 7489 23097 7523 23121
rect 7534 23097 7606 23131
rect 7489 23087 7606 23097
rect 7261 23063 7606 23087
rect 7274 23019 7474 23063
rect 7489 23053 7513 23063
rect 7489 23029 7523 23053
rect 7534 23029 7606 23063
rect 7489 23019 7606 23029
rect 7261 22995 7606 23019
rect 7274 22951 7474 22995
rect 7489 22985 7513 22995
rect 7489 22961 7523 22985
rect 7534 22961 7606 22995
rect 7489 22951 7606 22961
rect 7261 22927 7606 22951
rect 7274 22915 7474 22927
rect 7285 22903 7309 22915
rect 7489 22903 7513 22927
rect 7534 22915 7606 22927
rect 7836 22915 7892 23915
rect 7908 22915 7964 23915
rect 8266 23835 8466 23915
rect 8481 23845 8515 23869
rect 8526 23845 8598 23915
rect 8481 23835 8598 23845
rect 8253 23811 8598 23835
rect 8266 23767 8466 23811
rect 8481 23801 8505 23811
rect 8481 23777 8515 23801
rect 8526 23777 8598 23811
rect 8481 23767 8598 23777
rect 8253 23743 8598 23767
rect 8266 23699 8466 23743
rect 8481 23733 8505 23743
rect 8481 23709 8515 23733
rect 8526 23709 8598 23743
rect 8481 23699 8598 23709
rect 8253 23675 8598 23699
rect 8266 23631 8466 23675
rect 8481 23665 8505 23675
rect 8481 23641 8515 23665
rect 8526 23641 8598 23675
rect 8481 23631 8598 23641
rect 8253 23607 8598 23631
rect 8266 23563 8466 23607
rect 8481 23597 8505 23607
rect 8481 23573 8515 23597
rect 8526 23573 8598 23607
rect 8481 23563 8598 23573
rect 8253 23539 8598 23563
rect 8266 23495 8466 23539
rect 8481 23529 8505 23539
rect 8481 23505 8515 23529
rect 8526 23505 8598 23539
rect 8481 23495 8598 23505
rect 8253 23471 8598 23495
rect 8266 23427 8466 23471
rect 8481 23461 8505 23471
rect 8481 23437 8515 23461
rect 8526 23437 8598 23471
rect 8481 23427 8598 23437
rect 8253 23403 8598 23427
rect 8266 23359 8466 23403
rect 8481 23393 8505 23403
rect 8481 23369 8515 23393
rect 8526 23369 8598 23403
rect 8481 23359 8598 23369
rect 8253 23335 8598 23359
rect 8266 23291 8466 23335
rect 8481 23325 8505 23335
rect 8481 23301 8515 23325
rect 8526 23301 8598 23335
rect 8481 23291 8598 23301
rect 8253 23267 8598 23291
rect 8266 23223 8466 23267
rect 8481 23257 8505 23267
rect 8481 23233 8515 23257
rect 8526 23233 8598 23267
rect 8481 23223 8598 23233
rect 8253 23199 8598 23223
rect 8266 23155 8466 23199
rect 8481 23189 8505 23199
rect 8481 23165 8515 23189
rect 8526 23165 8598 23199
rect 8481 23155 8598 23165
rect 8253 23131 8598 23155
rect 8266 23087 8466 23131
rect 8481 23121 8505 23131
rect 8481 23097 8515 23121
rect 8526 23097 8598 23131
rect 8481 23087 8598 23097
rect 8253 23063 8598 23087
rect 8266 23019 8466 23063
rect 8481 23053 8505 23063
rect 8481 23029 8515 23053
rect 8526 23029 8598 23063
rect 8481 23019 8598 23029
rect 8253 22995 8598 23019
rect 8266 22951 8466 22995
rect 8481 22985 8505 22995
rect 8481 22961 8515 22985
rect 8526 22961 8598 22995
rect 8481 22951 8598 22961
rect 8253 22927 8598 22951
rect 8266 22915 8466 22927
rect 8277 22903 8301 22915
rect 8481 22903 8505 22927
rect 8526 22915 8598 22927
rect 8828 22915 8884 23915
rect 8900 22915 8956 23915
rect 9258 23835 9458 23915
rect 9473 23845 9507 23869
rect 9518 23845 9590 23915
rect 9473 23835 9590 23845
rect 9245 23811 9590 23835
rect 9258 23767 9458 23811
rect 9473 23801 9497 23811
rect 9473 23777 9507 23801
rect 9518 23777 9590 23811
rect 9473 23767 9590 23777
rect 9245 23743 9590 23767
rect 9258 23699 9458 23743
rect 9473 23733 9497 23743
rect 9473 23709 9507 23733
rect 9518 23709 9590 23743
rect 9473 23699 9590 23709
rect 9245 23675 9590 23699
rect 9258 23631 9458 23675
rect 9473 23665 9497 23675
rect 9473 23641 9507 23665
rect 9518 23641 9590 23675
rect 9473 23631 9590 23641
rect 9245 23607 9590 23631
rect 9258 23563 9458 23607
rect 9473 23597 9497 23607
rect 9473 23573 9507 23597
rect 9518 23573 9590 23607
rect 9473 23563 9590 23573
rect 9245 23539 9590 23563
rect 9258 23495 9458 23539
rect 9473 23529 9497 23539
rect 9473 23505 9507 23529
rect 9518 23505 9590 23539
rect 9473 23495 9590 23505
rect 9245 23471 9590 23495
rect 9258 23427 9458 23471
rect 9473 23461 9497 23471
rect 9473 23437 9507 23461
rect 9518 23437 9590 23471
rect 9473 23427 9590 23437
rect 9245 23403 9590 23427
rect 9258 23359 9458 23403
rect 9473 23393 9497 23403
rect 9473 23369 9507 23393
rect 9518 23369 9590 23403
rect 9473 23359 9590 23369
rect 9245 23335 9590 23359
rect 9258 23291 9458 23335
rect 9473 23325 9497 23335
rect 9473 23301 9507 23325
rect 9518 23301 9590 23335
rect 9473 23291 9590 23301
rect 9245 23267 9590 23291
rect 9258 23223 9458 23267
rect 9473 23257 9497 23267
rect 9473 23233 9507 23257
rect 9518 23233 9590 23267
rect 9473 23223 9590 23233
rect 9245 23199 9590 23223
rect 9258 23155 9458 23199
rect 9473 23189 9497 23199
rect 9473 23165 9507 23189
rect 9518 23165 9590 23199
rect 9473 23155 9590 23165
rect 9245 23131 9590 23155
rect 9258 23087 9458 23131
rect 9473 23121 9497 23131
rect 9473 23097 9507 23121
rect 9518 23097 9590 23131
rect 9473 23087 9590 23097
rect 9245 23063 9590 23087
rect 9258 23019 9458 23063
rect 9473 23053 9497 23063
rect 9473 23029 9507 23053
rect 9518 23029 9590 23063
rect 9473 23019 9590 23029
rect 9245 22995 9590 23019
rect 9258 22951 9458 22995
rect 9473 22985 9497 22995
rect 9473 22961 9507 22985
rect 9518 22961 9590 22995
rect 9473 22951 9590 22961
rect 9245 22927 9590 22951
rect 9258 22915 9458 22927
rect 9269 22903 9293 22915
rect 9473 22903 9497 22927
rect 9518 22915 9590 22927
rect 9820 22915 9876 23915
rect 9892 22915 9948 23915
rect 10250 23835 10450 23915
rect 10465 23845 10499 23869
rect 10510 23845 10582 23915
rect 10465 23835 10582 23845
rect 10237 23811 10582 23835
rect 10250 23767 10450 23811
rect 10465 23801 10489 23811
rect 10465 23777 10499 23801
rect 10510 23777 10582 23811
rect 10465 23767 10582 23777
rect 10237 23743 10582 23767
rect 10250 23699 10450 23743
rect 10465 23733 10489 23743
rect 10465 23709 10499 23733
rect 10510 23709 10582 23743
rect 10465 23699 10582 23709
rect 10237 23675 10582 23699
rect 10250 23631 10450 23675
rect 10465 23665 10489 23675
rect 10465 23641 10499 23665
rect 10510 23641 10582 23675
rect 10465 23631 10582 23641
rect 10237 23607 10582 23631
rect 10250 23563 10450 23607
rect 10465 23597 10489 23607
rect 10465 23573 10499 23597
rect 10510 23573 10582 23607
rect 10465 23563 10582 23573
rect 10237 23539 10582 23563
rect 10250 23495 10450 23539
rect 10465 23529 10489 23539
rect 10465 23505 10499 23529
rect 10510 23505 10582 23539
rect 10465 23495 10582 23505
rect 10237 23471 10582 23495
rect 10250 23427 10450 23471
rect 10465 23461 10489 23471
rect 10465 23437 10499 23461
rect 10510 23437 10582 23471
rect 10465 23427 10582 23437
rect 10237 23403 10582 23427
rect 10250 23359 10450 23403
rect 10465 23393 10489 23403
rect 10465 23369 10499 23393
rect 10510 23369 10582 23403
rect 10465 23359 10582 23369
rect 10237 23335 10582 23359
rect 10250 23291 10450 23335
rect 10465 23325 10489 23335
rect 10465 23301 10499 23325
rect 10510 23301 10582 23335
rect 10465 23291 10582 23301
rect 10237 23267 10582 23291
rect 10250 23223 10450 23267
rect 10465 23257 10489 23267
rect 10465 23233 10499 23257
rect 10510 23233 10582 23267
rect 10465 23223 10582 23233
rect 10237 23199 10582 23223
rect 10250 23155 10450 23199
rect 10465 23189 10489 23199
rect 10465 23165 10499 23189
rect 10510 23165 10582 23199
rect 10465 23155 10582 23165
rect 10237 23131 10582 23155
rect 10250 23087 10450 23131
rect 10465 23121 10489 23131
rect 10465 23097 10499 23121
rect 10510 23097 10582 23131
rect 10465 23087 10582 23097
rect 10237 23063 10582 23087
rect 10250 23019 10450 23063
rect 10465 23053 10489 23063
rect 10465 23029 10499 23053
rect 10510 23029 10582 23063
rect 10465 23019 10582 23029
rect 10237 22995 10582 23019
rect 10250 22951 10450 22995
rect 10465 22985 10489 22995
rect 10465 22961 10499 22985
rect 10510 22961 10582 22995
rect 10465 22951 10582 22961
rect 10237 22927 10582 22951
rect 10250 22915 10450 22927
rect 10261 22903 10285 22915
rect 10465 22903 10489 22927
rect 10510 22915 10582 22927
rect 10812 22915 10868 23915
rect 10884 22915 10940 23915
rect 11242 23835 11442 23915
rect 11457 23845 11491 23869
rect 11502 23845 11574 23915
rect 11457 23835 11574 23845
rect 11229 23811 11574 23835
rect 11242 23767 11442 23811
rect 11457 23801 11481 23811
rect 11457 23777 11491 23801
rect 11502 23777 11574 23811
rect 11457 23767 11574 23777
rect 11229 23743 11574 23767
rect 11242 23699 11442 23743
rect 11457 23733 11481 23743
rect 11457 23709 11491 23733
rect 11502 23709 11574 23743
rect 11457 23699 11574 23709
rect 11229 23675 11574 23699
rect 11242 23631 11442 23675
rect 11457 23665 11481 23675
rect 11457 23641 11491 23665
rect 11502 23641 11574 23675
rect 11457 23631 11574 23641
rect 11229 23607 11574 23631
rect 11242 23563 11442 23607
rect 11457 23597 11481 23607
rect 11457 23573 11491 23597
rect 11502 23573 11574 23607
rect 11457 23563 11574 23573
rect 11229 23539 11574 23563
rect 11242 23495 11442 23539
rect 11457 23529 11481 23539
rect 11457 23505 11491 23529
rect 11502 23505 11574 23539
rect 11457 23495 11574 23505
rect 11229 23471 11574 23495
rect 11242 23427 11442 23471
rect 11457 23461 11481 23471
rect 11457 23437 11491 23461
rect 11502 23437 11574 23471
rect 11457 23427 11574 23437
rect 11229 23403 11574 23427
rect 11242 23359 11442 23403
rect 11457 23393 11481 23403
rect 11457 23369 11491 23393
rect 11502 23369 11574 23403
rect 11457 23359 11574 23369
rect 11229 23335 11574 23359
rect 11242 23291 11442 23335
rect 11457 23325 11481 23335
rect 11457 23301 11491 23325
rect 11502 23301 11574 23335
rect 11457 23291 11574 23301
rect 11229 23267 11574 23291
rect 11242 23223 11442 23267
rect 11457 23257 11481 23267
rect 11457 23233 11491 23257
rect 11502 23233 11574 23267
rect 11457 23223 11574 23233
rect 11229 23199 11574 23223
rect 11242 23155 11442 23199
rect 11457 23189 11481 23199
rect 11457 23165 11491 23189
rect 11502 23165 11574 23199
rect 11457 23155 11574 23165
rect 11229 23131 11574 23155
rect 11242 23087 11442 23131
rect 11457 23121 11481 23131
rect 11457 23097 11491 23121
rect 11502 23097 11574 23131
rect 11457 23087 11574 23097
rect 11229 23063 11574 23087
rect 11242 23019 11442 23063
rect 11457 23053 11481 23063
rect 11457 23029 11491 23053
rect 11502 23029 11574 23063
rect 11457 23019 11574 23029
rect 11229 22995 11574 23019
rect 11242 22951 11442 22995
rect 11457 22985 11481 22995
rect 11457 22961 11491 22985
rect 11502 22961 11574 22995
rect 11457 22951 11574 22961
rect 11229 22927 11574 22951
rect 11242 22915 11442 22927
rect 11253 22903 11277 22915
rect 11457 22903 11481 22927
rect 11502 22915 11574 22927
rect 11804 22915 11860 23915
rect 11876 22915 11932 23915
rect 12234 23835 12434 23915
rect 12449 23845 12483 23869
rect 12494 23845 12566 23915
rect 12449 23835 12566 23845
rect 12221 23811 12566 23835
rect 12234 23767 12434 23811
rect 12449 23801 12473 23811
rect 12449 23777 12483 23801
rect 12494 23777 12566 23811
rect 12449 23767 12566 23777
rect 12221 23743 12566 23767
rect 12234 23699 12434 23743
rect 12449 23733 12473 23743
rect 12449 23709 12483 23733
rect 12494 23709 12566 23743
rect 12449 23699 12566 23709
rect 12221 23675 12566 23699
rect 12234 23631 12434 23675
rect 12449 23665 12473 23675
rect 12449 23641 12483 23665
rect 12494 23641 12566 23675
rect 12449 23631 12566 23641
rect 12221 23607 12566 23631
rect 12234 23563 12434 23607
rect 12449 23597 12473 23607
rect 12449 23573 12483 23597
rect 12494 23573 12566 23607
rect 12449 23563 12566 23573
rect 12221 23539 12566 23563
rect 12234 23495 12434 23539
rect 12449 23529 12473 23539
rect 12449 23505 12483 23529
rect 12494 23505 12566 23539
rect 12449 23495 12566 23505
rect 12221 23471 12566 23495
rect 12234 23427 12434 23471
rect 12449 23461 12473 23471
rect 12449 23437 12483 23461
rect 12494 23437 12566 23471
rect 12449 23427 12566 23437
rect 12221 23403 12566 23427
rect 12234 23359 12434 23403
rect 12449 23393 12473 23403
rect 12449 23369 12483 23393
rect 12494 23369 12566 23403
rect 12449 23359 12566 23369
rect 12221 23335 12566 23359
rect 12234 23291 12434 23335
rect 12449 23325 12473 23335
rect 12449 23301 12483 23325
rect 12494 23301 12566 23335
rect 12449 23291 12566 23301
rect 12221 23267 12566 23291
rect 12234 23223 12434 23267
rect 12449 23257 12473 23267
rect 12449 23233 12483 23257
rect 12494 23233 12566 23267
rect 12449 23223 12566 23233
rect 12221 23199 12566 23223
rect 12234 23155 12434 23199
rect 12449 23189 12473 23199
rect 12449 23165 12483 23189
rect 12494 23165 12566 23199
rect 12449 23155 12566 23165
rect 12221 23131 12566 23155
rect 12234 23087 12434 23131
rect 12449 23121 12473 23131
rect 12449 23097 12483 23121
rect 12494 23097 12566 23131
rect 12449 23087 12566 23097
rect 12221 23063 12566 23087
rect 12234 23019 12434 23063
rect 12449 23053 12473 23063
rect 12449 23029 12483 23053
rect 12494 23029 12566 23063
rect 12449 23019 12566 23029
rect 12221 22995 12566 23019
rect 12234 22951 12434 22995
rect 12449 22985 12473 22995
rect 12449 22961 12483 22985
rect 12494 22961 12566 22995
rect 12449 22951 12566 22961
rect 12221 22927 12566 22951
rect 12234 22915 12434 22927
rect 12245 22903 12269 22915
rect 12449 22903 12473 22927
rect 12494 22915 12566 22927
rect 12796 22915 12852 23915
rect 12868 22915 12924 23915
rect 13226 23835 13426 23915
rect 13441 23845 13475 23869
rect 13486 23845 13558 23915
rect 13441 23835 13558 23845
rect 13213 23811 13558 23835
rect 13226 23767 13426 23811
rect 13441 23801 13465 23811
rect 13441 23777 13475 23801
rect 13486 23777 13558 23811
rect 13441 23767 13558 23777
rect 13213 23743 13558 23767
rect 13226 23699 13426 23743
rect 13441 23733 13465 23743
rect 13441 23709 13475 23733
rect 13486 23709 13558 23743
rect 13441 23699 13558 23709
rect 13213 23675 13558 23699
rect 13226 23631 13426 23675
rect 13441 23665 13465 23675
rect 13441 23641 13475 23665
rect 13486 23641 13558 23675
rect 13441 23631 13558 23641
rect 13213 23607 13558 23631
rect 13226 23563 13426 23607
rect 13441 23597 13465 23607
rect 13441 23573 13475 23597
rect 13486 23573 13558 23607
rect 13441 23563 13558 23573
rect 13213 23539 13558 23563
rect 13226 23495 13426 23539
rect 13441 23529 13465 23539
rect 13441 23505 13475 23529
rect 13486 23505 13558 23539
rect 13441 23495 13558 23505
rect 13213 23471 13558 23495
rect 13226 23427 13426 23471
rect 13441 23461 13465 23471
rect 13441 23437 13475 23461
rect 13486 23437 13558 23471
rect 13441 23427 13558 23437
rect 13213 23403 13558 23427
rect 13226 23359 13426 23403
rect 13441 23393 13465 23403
rect 13441 23369 13475 23393
rect 13486 23369 13558 23403
rect 13441 23359 13558 23369
rect 13213 23335 13558 23359
rect 13226 23291 13426 23335
rect 13441 23325 13465 23335
rect 13441 23301 13475 23325
rect 13486 23301 13558 23335
rect 13441 23291 13558 23301
rect 13213 23267 13558 23291
rect 13226 23223 13426 23267
rect 13441 23257 13465 23267
rect 13441 23233 13475 23257
rect 13486 23233 13558 23267
rect 13441 23223 13558 23233
rect 13213 23199 13558 23223
rect 13226 23155 13426 23199
rect 13441 23189 13465 23199
rect 13441 23165 13475 23189
rect 13486 23165 13558 23199
rect 13441 23155 13558 23165
rect 13213 23131 13558 23155
rect 13226 23087 13426 23131
rect 13441 23121 13465 23131
rect 13441 23097 13475 23121
rect 13486 23097 13558 23131
rect 13441 23087 13558 23097
rect 13213 23063 13558 23087
rect 13226 23019 13426 23063
rect 13441 23053 13465 23063
rect 13441 23029 13475 23053
rect 13486 23029 13558 23063
rect 13441 23019 13558 23029
rect 13213 22995 13558 23019
rect 13226 22951 13426 22995
rect 13441 22985 13465 22995
rect 13441 22961 13475 22985
rect 13486 22961 13558 22995
rect 13441 22951 13558 22961
rect 13213 22927 13558 22951
rect 13226 22915 13426 22927
rect 13237 22903 13261 22915
rect 13441 22903 13465 22927
rect 13486 22915 13558 22927
rect 13788 22915 13844 23915
rect 13860 22915 13916 23915
rect 14218 23835 14418 23915
rect 14433 23845 14467 23869
rect 14478 23845 14550 23915
rect 14433 23835 14550 23845
rect 14205 23811 14550 23835
rect 14218 23767 14418 23811
rect 14433 23801 14457 23811
rect 14433 23777 14467 23801
rect 14478 23777 14550 23811
rect 14433 23767 14550 23777
rect 14205 23743 14550 23767
rect 14218 23699 14418 23743
rect 14433 23733 14457 23743
rect 14433 23709 14467 23733
rect 14478 23709 14550 23743
rect 14433 23699 14550 23709
rect 14205 23675 14550 23699
rect 14218 23631 14418 23675
rect 14433 23665 14457 23675
rect 14433 23641 14467 23665
rect 14478 23641 14550 23675
rect 14433 23631 14550 23641
rect 14205 23607 14550 23631
rect 14218 23563 14418 23607
rect 14433 23597 14457 23607
rect 14433 23573 14467 23597
rect 14478 23573 14550 23607
rect 14433 23563 14550 23573
rect 14205 23539 14550 23563
rect 14218 23495 14418 23539
rect 14433 23529 14457 23539
rect 14433 23505 14467 23529
rect 14478 23505 14550 23539
rect 14433 23495 14550 23505
rect 14205 23471 14550 23495
rect 14218 23427 14418 23471
rect 14433 23461 14457 23471
rect 14433 23437 14467 23461
rect 14478 23437 14550 23471
rect 14433 23427 14550 23437
rect 14205 23403 14550 23427
rect 14218 23359 14418 23403
rect 14433 23393 14457 23403
rect 14433 23369 14467 23393
rect 14478 23369 14550 23403
rect 14433 23359 14550 23369
rect 14205 23335 14550 23359
rect 14218 23291 14418 23335
rect 14433 23325 14457 23335
rect 14433 23301 14467 23325
rect 14478 23301 14550 23335
rect 14433 23291 14550 23301
rect 14205 23267 14550 23291
rect 14218 23223 14418 23267
rect 14433 23257 14457 23267
rect 14433 23233 14467 23257
rect 14478 23233 14550 23267
rect 14433 23223 14550 23233
rect 14205 23199 14550 23223
rect 14218 23155 14418 23199
rect 14433 23189 14457 23199
rect 14433 23165 14467 23189
rect 14478 23165 14550 23199
rect 14433 23155 14550 23165
rect 14205 23131 14550 23155
rect 14218 23087 14418 23131
rect 14433 23121 14457 23131
rect 14433 23097 14467 23121
rect 14478 23097 14550 23131
rect 14433 23087 14550 23097
rect 14205 23063 14550 23087
rect 14218 23019 14418 23063
rect 14433 23053 14457 23063
rect 14433 23029 14467 23053
rect 14478 23029 14550 23063
rect 14433 23019 14550 23029
rect 14205 22995 14550 23019
rect 14218 22951 14418 22995
rect 14433 22985 14457 22995
rect 14433 22961 14467 22985
rect 14478 22961 14550 22995
rect 14433 22951 14550 22961
rect 14205 22927 14550 22951
rect 14218 22915 14418 22927
rect 14229 22903 14253 22915
rect 14433 22903 14457 22927
rect 14478 22915 14550 22927
rect 14739 22915 14811 23915
rect 14877 22915 14894 23915
rect 15064 22915 15097 23915
rect 15220 23723 15288 23749
rect 15220 23689 15254 23715
rect 2325 22315 2359 22327
rect 1623 21315 1673 22315
rect 1884 21315 1940 22315
rect 1956 21315 2012 22315
rect 2314 22293 2514 22315
rect 2529 22303 2563 22327
rect 3317 22315 3351 22327
rect 2574 22303 2646 22315
rect 2529 22293 2646 22303
rect 2301 22269 2646 22293
rect 2314 22225 2514 22269
rect 2529 22259 2553 22269
rect 2529 22235 2563 22259
rect 2574 22235 2646 22269
rect 2529 22225 2646 22235
rect 2301 22201 2646 22225
rect 2314 22157 2514 22201
rect 2529 22191 2553 22201
rect 2529 22167 2563 22191
rect 2574 22167 2646 22201
rect 2529 22157 2646 22167
rect 2301 22133 2646 22157
rect 2314 22089 2514 22133
rect 2529 22123 2553 22133
rect 2529 22099 2563 22123
rect 2574 22099 2646 22133
rect 2529 22089 2646 22099
rect 2301 22065 2646 22089
rect 2314 22021 2514 22065
rect 2529 22055 2553 22065
rect 2529 22031 2563 22055
rect 2574 22031 2646 22065
rect 2529 22021 2646 22031
rect 2301 21997 2646 22021
rect 2314 21953 2514 21997
rect 2529 21987 2553 21997
rect 2529 21963 2563 21987
rect 2574 21963 2646 21997
rect 2529 21953 2646 21963
rect 2301 21929 2646 21953
rect 2314 21885 2514 21929
rect 2529 21919 2553 21929
rect 2529 21895 2563 21919
rect 2574 21895 2646 21929
rect 2529 21885 2646 21895
rect 2301 21861 2646 21885
rect 2314 21817 2514 21861
rect 2529 21851 2553 21861
rect 2529 21827 2563 21851
rect 2574 21827 2646 21861
rect 2529 21817 2646 21827
rect 2301 21793 2646 21817
rect 2314 21749 2514 21793
rect 2529 21783 2553 21793
rect 2529 21759 2563 21783
rect 2574 21759 2646 21793
rect 2529 21749 2646 21759
rect 2301 21725 2646 21749
rect 2314 21681 2514 21725
rect 2529 21715 2553 21725
rect 2529 21691 2563 21715
rect 2574 21691 2646 21725
rect 2529 21681 2646 21691
rect 2301 21657 2646 21681
rect 2314 21613 2514 21657
rect 2529 21647 2553 21657
rect 2529 21623 2563 21647
rect 2574 21623 2646 21657
rect 2529 21613 2646 21623
rect 2301 21589 2646 21613
rect 2314 21545 2514 21589
rect 2529 21579 2553 21589
rect 2529 21555 2563 21579
rect 2574 21555 2646 21589
rect 2529 21545 2646 21555
rect 2301 21521 2646 21545
rect 2314 21477 2514 21521
rect 2529 21511 2553 21521
rect 2529 21487 2563 21511
rect 2574 21487 2646 21521
rect 2529 21477 2646 21487
rect 2301 21453 2646 21477
rect 2314 21409 2514 21453
rect 2529 21443 2553 21453
rect 2529 21419 2563 21443
rect 2574 21419 2646 21453
rect 2529 21409 2646 21419
rect 2301 21385 2646 21409
rect 2314 21315 2514 21385
rect 2529 21361 2553 21385
rect 2574 21315 2646 21385
rect 2876 21315 2932 22315
rect 2948 21315 3004 22315
rect 3306 22293 3506 22315
rect 3521 22303 3555 22327
rect 4309 22315 4343 22327
rect 3566 22303 3638 22315
rect 3521 22293 3638 22303
rect 3293 22269 3638 22293
rect 3306 22225 3506 22269
rect 3521 22259 3545 22269
rect 3521 22235 3555 22259
rect 3566 22235 3638 22269
rect 3521 22225 3638 22235
rect 3293 22201 3638 22225
rect 3306 22157 3506 22201
rect 3521 22191 3545 22201
rect 3521 22167 3555 22191
rect 3566 22167 3638 22201
rect 3521 22157 3638 22167
rect 3293 22133 3638 22157
rect 3306 22089 3506 22133
rect 3521 22123 3545 22133
rect 3521 22099 3555 22123
rect 3566 22099 3638 22133
rect 3521 22089 3638 22099
rect 3293 22065 3638 22089
rect 3306 22021 3506 22065
rect 3521 22055 3545 22065
rect 3521 22031 3555 22055
rect 3566 22031 3638 22065
rect 3521 22021 3638 22031
rect 3293 21997 3638 22021
rect 3306 21953 3506 21997
rect 3521 21987 3545 21997
rect 3521 21963 3555 21987
rect 3566 21963 3638 21997
rect 3521 21953 3638 21963
rect 3293 21929 3638 21953
rect 3306 21885 3506 21929
rect 3521 21919 3545 21929
rect 3521 21895 3555 21919
rect 3566 21895 3638 21929
rect 3521 21885 3638 21895
rect 3293 21861 3638 21885
rect 3306 21817 3506 21861
rect 3521 21851 3545 21861
rect 3521 21827 3555 21851
rect 3566 21827 3638 21861
rect 3521 21817 3638 21827
rect 3293 21793 3638 21817
rect 3306 21749 3506 21793
rect 3521 21783 3545 21793
rect 3521 21759 3555 21783
rect 3566 21759 3638 21793
rect 3521 21749 3638 21759
rect 3293 21725 3638 21749
rect 3306 21681 3506 21725
rect 3521 21715 3545 21725
rect 3521 21691 3555 21715
rect 3566 21691 3638 21725
rect 3521 21681 3638 21691
rect 3293 21657 3638 21681
rect 3306 21613 3506 21657
rect 3521 21647 3545 21657
rect 3521 21623 3555 21647
rect 3566 21623 3638 21657
rect 3521 21613 3638 21623
rect 3293 21589 3638 21613
rect 3306 21545 3506 21589
rect 3521 21579 3545 21589
rect 3521 21555 3555 21579
rect 3566 21555 3638 21589
rect 3521 21545 3638 21555
rect 3293 21521 3638 21545
rect 3306 21477 3506 21521
rect 3521 21511 3545 21521
rect 3521 21487 3555 21511
rect 3566 21487 3638 21521
rect 3521 21477 3638 21487
rect 3293 21453 3638 21477
rect 3306 21409 3506 21453
rect 3521 21443 3545 21453
rect 3521 21419 3555 21443
rect 3566 21419 3638 21453
rect 3521 21409 3638 21419
rect 3293 21385 3638 21409
rect 3306 21315 3506 21385
rect 3521 21361 3545 21385
rect 3566 21315 3638 21385
rect 3868 21315 3924 22315
rect 3940 21315 3996 22315
rect 4298 22293 4498 22315
rect 4513 22303 4547 22327
rect 5301 22315 5335 22327
rect 4558 22303 4630 22315
rect 4513 22293 4630 22303
rect 4285 22269 4630 22293
rect 4298 22225 4498 22269
rect 4513 22259 4537 22269
rect 4513 22235 4547 22259
rect 4558 22235 4630 22269
rect 4513 22225 4630 22235
rect 4285 22201 4630 22225
rect 4298 22157 4498 22201
rect 4513 22191 4537 22201
rect 4513 22167 4547 22191
rect 4558 22167 4630 22201
rect 4513 22157 4630 22167
rect 4285 22133 4630 22157
rect 4298 22089 4498 22133
rect 4513 22123 4537 22133
rect 4513 22099 4547 22123
rect 4558 22099 4630 22133
rect 4513 22089 4630 22099
rect 4285 22065 4630 22089
rect 4298 22021 4498 22065
rect 4513 22055 4537 22065
rect 4513 22031 4547 22055
rect 4558 22031 4630 22065
rect 4513 22021 4630 22031
rect 4285 21997 4630 22021
rect 4298 21953 4498 21997
rect 4513 21987 4537 21997
rect 4513 21963 4547 21987
rect 4558 21963 4630 21997
rect 4513 21953 4630 21963
rect 4285 21929 4630 21953
rect 4298 21885 4498 21929
rect 4513 21919 4537 21929
rect 4513 21895 4547 21919
rect 4558 21895 4630 21929
rect 4513 21885 4630 21895
rect 4285 21861 4630 21885
rect 4298 21817 4498 21861
rect 4513 21851 4537 21861
rect 4513 21827 4547 21851
rect 4558 21827 4630 21861
rect 4513 21817 4630 21827
rect 4285 21793 4630 21817
rect 4298 21749 4498 21793
rect 4513 21783 4537 21793
rect 4513 21759 4547 21783
rect 4558 21759 4630 21793
rect 4513 21749 4630 21759
rect 4285 21725 4630 21749
rect 4298 21681 4498 21725
rect 4513 21715 4537 21725
rect 4513 21691 4547 21715
rect 4558 21691 4630 21725
rect 4513 21681 4630 21691
rect 4285 21657 4630 21681
rect 4298 21613 4498 21657
rect 4513 21647 4537 21657
rect 4513 21623 4547 21647
rect 4558 21623 4630 21657
rect 4513 21613 4630 21623
rect 4285 21589 4630 21613
rect 4298 21545 4498 21589
rect 4513 21579 4537 21589
rect 4513 21555 4547 21579
rect 4558 21555 4630 21589
rect 4513 21545 4630 21555
rect 4285 21521 4630 21545
rect 4298 21477 4498 21521
rect 4513 21511 4537 21521
rect 4513 21487 4547 21511
rect 4558 21487 4630 21521
rect 4513 21477 4630 21487
rect 4285 21453 4630 21477
rect 4298 21409 4498 21453
rect 4513 21443 4537 21453
rect 4513 21419 4547 21443
rect 4558 21419 4630 21453
rect 4513 21409 4630 21419
rect 4285 21385 4630 21409
rect 4298 21315 4498 21385
rect 4513 21361 4537 21385
rect 4558 21315 4630 21385
rect 4860 21315 4916 22315
rect 4932 21315 4988 22315
rect 5290 22293 5490 22315
rect 5505 22303 5539 22327
rect 6293 22315 6327 22327
rect 5550 22303 5622 22315
rect 5505 22293 5622 22303
rect 5277 22269 5622 22293
rect 5290 22225 5490 22269
rect 5505 22259 5529 22269
rect 5505 22235 5539 22259
rect 5550 22235 5622 22269
rect 5505 22225 5622 22235
rect 5277 22201 5622 22225
rect 5290 22157 5490 22201
rect 5505 22191 5529 22201
rect 5505 22167 5539 22191
rect 5550 22167 5622 22201
rect 5505 22157 5622 22167
rect 5277 22133 5622 22157
rect 5290 22089 5490 22133
rect 5505 22123 5529 22133
rect 5505 22099 5539 22123
rect 5550 22099 5622 22133
rect 5505 22089 5622 22099
rect 5277 22065 5622 22089
rect 5290 22021 5490 22065
rect 5505 22055 5529 22065
rect 5505 22031 5539 22055
rect 5550 22031 5622 22065
rect 5505 22021 5622 22031
rect 5277 21997 5622 22021
rect 5290 21953 5490 21997
rect 5505 21987 5529 21997
rect 5505 21963 5539 21987
rect 5550 21963 5622 21997
rect 5505 21953 5622 21963
rect 5277 21929 5622 21953
rect 5290 21885 5490 21929
rect 5505 21919 5529 21929
rect 5505 21895 5539 21919
rect 5550 21895 5622 21929
rect 5505 21885 5622 21895
rect 5277 21861 5622 21885
rect 5290 21817 5490 21861
rect 5505 21851 5529 21861
rect 5505 21827 5539 21851
rect 5550 21827 5622 21861
rect 5505 21817 5622 21827
rect 5277 21793 5622 21817
rect 5290 21749 5490 21793
rect 5505 21783 5529 21793
rect 5505 21759 5539 21783
rect 5550 21759 5622 21793
rect 5505 21749 5622 21759
rect 5277 21725 5622 21749
rect 5290 21681 5490 21725
rect 5505 21715 5529 21725
rect 5505 21691 5539 21715
rect 5550 21691 5622 21725
rect 5505 21681 5622 21691
rect 5277 21657 5622 21681
rect 5290 21613 5490 21657
rect 5505 21647 5529 21657
rect 5505 21623 5539 21647
rect 5550 21623 5622 21657
rect 5505 21613 5622 21623
rect 5277 21589 5622 21613
rect 5290 21545 5490 21589
rect 5505 21579 5529 21589
rect 5505 21555 5539 21579
rect 5550 21555 5622 21589
rect 5505 21545 5622 21555
rect 5277 21521 5622 21545
rect 5290 21477 5490 21521
rect 5505 21511 5529 21521
rect 5505 21487 5539 21511
rect 5550 21487 5622 21521
rect 5505 21477 5622 21487
rect 5277 21453 5622 21477
rect 5290 21409 5490 21453
rect 5505 21443 5529 21453
rect 5505 21419 5539 21443
rect 5550 21419 5622 21453
rect 5505 21409 5622 21419
rect 5277 21385 5622 21409
rect 5290 21315 5490 21385
rect 5505 21361 5529 21385
rect 5550 21315 5622 21385
rect 5852 21315 5908 22315
rect 5924 21315 5980 22315
rect 6282 22293 6482 22315
rect 6497 22303 6531 22327
rect 7285 22315 7319 22327
rect 6542 22303 6614 22315
rect 6497 22293 6614 22303
rect 6269 22269 6614 22293
rect 6282 22225 6482 22269
rect 6497 22259 6521 22269
rect 6497 22235 6531 22259
rect 6542 22235 6614 22269
rect 6497 22225 6614 22235
rect 6269 22201 6614 22225
rect 6282 22157 6482 22201
rect 6497 22191 6521 22201
rect 6497 22167 6531 22191
rect 6542 22167 6614 22201
rect 6497 22157 6614 22167
rect 6269 22133 6614 22157
rect 6282 22089 6482 22133
rect 6497 22123 6521 22133
rect 6497 22099 6531 22123
rect 6542 22099 6614 22133
rect 6497 22089 6614 22099
rect 6269 22065 6614 22089
rect 6282 22021 6482 22065
rect 6497 22055 6521 22065
rect 6497 22031 6531 22055
rect 6542 22031 6614 22065
rect 6497 22021 6614 22031
rect 6269 21997 6614 22021
rect 6282 21953 6482 21997
rect 6497 21987 6521 21997
rect 6497 21963 6531 21987
rect 6542 21963 6614 21997
rect 6497 21953 6614 21963
rect 6269 21929 6614 21953
rect 6282 21885 6482 21929
rect 6497 21919 6521 21929
rect 6497 21895 6531 21919
rect 6542 21895 6614 21929
rect 6497 21885 6614 21895
rect 6269 21861 6614 21885
rect 6282 21817 6482 21861
rect 6497 21851 6521 21861
rect 6497 21827 6531 21851
rect 6542 21827 6614 21861
rect 6497 21817 6614 21827
rect 6269 21793 6614 21817
rect 6282 21749 6482 21793
rect 6497 21783 6521 21793
rect 6497 21759 6531 21783
rect 6542 21759 6614 21793
rect 6497 21749 6614 21759
rect 6269 21725 6614 21749
rect 6282 21681 6482 21725
rect 6497 21715 6521 21725
rect 6497 21691 6531 21715
rect 6542 21691 6614 21725
rect 6497 21681 6614 21691
rect 6269 21657 6614 21681
rect 6282 21613 6482 21657
rect 6497 21647 6521 21657
rect 6497 21623 6531 21647
rect 6542 21623 6614 21657
rect 6497 21613 6614 21623
rect 6269 21589 6614 21613
rect 6282 21545 6482 21589
rect 6497 21579 6521 21589
rect 6497 21555 6531 21579
rect 6542 21555 6614 21589
rect 6497 21545 6614 21555
rect 6269 21521 6614 21545
rect 6282 21477 6482 21521
rect 6497 21511 6521 21521
rect 6497 21487 6531 21511
rect 6542 21487 6614 21521
rect 6497 21477 6614 21487
rect 6269 21453 6614 21477
rect 6282 21409 6482 21453
rect 6497 21443 6521 21453
rect 6497 21419 6531 21443
rect 6542 21419 6614 21453
rect 6497 21409 6614 21419
rect 6269 21385 6614 21409
rect 6282 21315 6482 21385
rect 6497 21361 6521 21385
rect 6542 21315 6614 21385
rect 6844 21315 6900 22315
rect 6916 21315 6972 22315
rect 7274 22293 7474 22315
rect 7489 22303 7523 22327
rect 8277 22315 8311 22327
rect 7534 22303 7606 22315
rect 7489 22293 7606 22303
rect 7261 22269 7606 22293
rect 7274 22225 7474 22269
rect 7489 22259 7513 22269
rect 7489 22235 7523 22259
rect 7534 22235 7606 22269
rect 7489 22225 7606 22235
rect 7261 22201 7606 22225
rect 7274 22157 7474 22201
rect 7489 22191 7513 22201
rect 7489 22167 7523 22191
rect 7534 22167 7606 22201
rect 7489 22157 7606 22167
rect 7261 22133 7606 22157
rect 7274 22089 7474 22133
rect 7489 22123 7513 22133
rect 7489 22099 7523 22123
rect 7534 22099 7606 22133
rect 7489 22089 7606 22099
rect 7261 22065 7606 22089
rect 7274 22021 7474 22065
rect 7489 22055 7513 22065
rect 7489 22031 7523 22055
rect 7534 22031 7606 22065
rect 7489 22021 7606 22031
rect 7261 21997 7606 22021
rect 7274 21953 7474 21997
rect 7489 21987 7513 21997
rect 7489 21963 7523 21987
rect 7534 21963 7606 21997
rect 7489 21953 7606 21963
rect 7261 21929 7606 21953
rect 7274 21885 7474 21929
rect 7489 21919 7513 21929
rect 7489 21895 7523 21919
rect 7534 21895 7606 21929
rect 7489 21885 7606 21895
rect 7261 21861 7606 21885
rect 7274 21817 7474 21861
rect 7489 21851 7513 21861
rect 7489 21827 7523 21851
rect 7534 21827 7606 21861
rect 7489 21817 7606 21827
rect 7261 21793 7606 21817
rect 7274 21749 7474 21793
rect 7489 21783 7513 21793
rect 7489 21759 7523 21783
rect 7534 21759 7606 21793
rect 7489 21749 7606 21759
rect 7261 21725 7606 21749
rect 7274 21681 7474 21725
rect 7489 21715 7513 21725
rect 7489 21691 7523 21715
rect 7534 21691 7606 21725
rect 7489 21681 7606 21691
rect 7261 21657 7606 21681
rect 7274 21613 7474 21657
rect 7489 21647 7513 21657
rect 7489 21623 7523 21647
rect 7534 21623 7606 21657
rect 7489 21613 7606 21623
rect 7261 21589 7606 21613
rect 7274 21545 7474 21589
rect 7489 21579 7513 21589
rect 7489 21555 7523 21579
rect 7534 21555 7606 21589
rect 7489 21545 7606 21555
rect 7261 21521 7606 21545
rect 7274 21477 7474 21521
rect 7489 21511 7513 21521
rect 7489 21487 7523 21511
rect 7534 21487 7606 21521
rect 7489 21477 7606 21487
rect 7261 21453 7606 21477
rect 7274 21409 7474 21453
rect 7489 21443 7513 21453
rect 7489 21419 7523 21443
rect 7534 21419 7606 21453
rect 7489 21409 7606 21419
rect 7261 21385 7606 21409
rect 7274 21315 7474 21385
rect 7489 21361 7513 21385
rect 7534 21315 7606 21385
rect 7836 21315 7892 22315
rect 7908 21315 7964 22315
rect 8266 22293 8466 22315
rect 8481 22303 8515 22327
rect 9269 22315 9303 22327
rect 8526 22303 8598 22315
rect 8481 22293 8598 22303
rect 8253 22269 8598 22293
rect 8266 22225 8466 22269
rect 8481 22259 8505 22269
rect 8481 22235 8515 22259
rect 8526 22235 8598 22269
rect 8481 22225 8598 22235
rect 8253 22201 8598 22225
rect 8266 22157 8466 22201
rect 8481 22191 8505 22201
rect 8481 22167 8515 22191
rect 8526 22167 8598 22201
rect 8481 22157 8598 22167
rect 8253 22133 8598 22157
rect 8266 22089 8466 22133
rect 8481 22123 8505 22133
rect 8481 22099 8515 22123
rect 8526 22099 8598 22133
rect 8481 22089 8598 22099
rect 8253 22065 8598 22089
rect 8266 22021 8466 22065
rect 8481 22055 8505 22065
rect 8481 22031 8515 22055
rect 8526 22031 8598 22065
rect 8481 22021 8598 22031
rect 8253 21997 8598 22021
rect 8266 21953 8466 21997
rect 8481 21987 8505 21997
rect 8481 21963 8515 21987
rect 8526 21963 8598 21997
rect 8481 21953 8598 21963
rect 8253 21929 8598 21953
rect 8266 21885 8466 21929
rect 8481 21919 8505 21929
rect 8481 21895 8515 21919
rect 8526 21895 8598 21929
rect 8481 21885 8598 21895
rect 8253 21861 8598 21885
rect 8266 21817 8466 21861
rect 8481 21851 8505 21861
rect 8481 21827 8515 21851
rect 8526 21827 8598 21861
rect 8481 21817 8598 21827
rect 8253 21793 8598 21817
rect 8266 21749 8466 21793
rect 8481 21783 8505 21793
rect 8481 21759 8515 21783
rect 8526 21759 8598 21793
rect 8481 21749 8598 21759
rect 8253 21725 8598 21749
rect 8266 21681 8466 21725
rect 8481 21715 8505 21725
rect 8481 21691 8515 21715
rect 8526 21691 8598 21725
rect 8481 21681 8598 21691
rect 8253 21657 8598 21681
rect 8266 21613 8466 21657
rect 8481 21647 8505 21657
rect 8481 21623 8515 21647
rect 8526 21623 8598 21657
rect 8481 21613 8598 21623
rect 8253 21589 8598 21613
rect 8266 21545 8466 21589
rect 8481 21579 8505 21589
rect 8481 21555 8515 21579
rect 8526 21555 8598 21589
rect 8481 21545 8598 21555
rect 8253 21521 8598 21545
rect 8266 21477 8466 21521
rect 8481 21511 8505 21521
rect 8481 21487 8515 21511
rect 8526 21487 8598 21521
rect 8481 21477 8598 21487
rect 8253 21453 8598 21477
rect 8266 21409 8466 21453
rect 8481 21443 8505 21453
rect 8481 21419 8515 21443
rect 8526 21419 8598 21453
rect 8481 21409 8598 21419
rect 8253 21385 8598 21409
rect 8266 21315 8466 21385
rect 8481 21361 8505 21385
rect 8526 21315 8598 21385
rect 8828 21315 8884 22315
rect 8900 21315 8956 22315
rect 9258 22293 9458 22315
rect 9473 22303 9507 22327
rect 10261 22315 10295 22327
rect 9518 22303 9590 22315
rect 9473 22293 9590 22303
rect 9245 22269 9590 22293
rect 9258 22225 9458 22269
rect 9473 22259 9497 22269
rect 9473 22235 9507 22259
rect 9518 22235 9590 22269
rect 9473 22225 9590 22235
rect 9245 22201 9590 22225
rect 9258 22157 9458 22201
rect 9473 22191 9497 22201
rect 9473 22167 9507 22191
rect 9518 22167 9590 22201
rect 9473 22157 9590 22167
rect 9245 22133 9590 22157
rect 9258 22089 9458 22133
rect 9473 22123 9497 22133
rect 9473 22099 9507 22123
rect 9518 22099 9590 22133
rect 9473 22089 9590 22099
rect 9245 22065 9590 22089
rect 9258 22021 9458 22065
rect 9473 22055 9497 22065
rect 9473 22031 9507 22055
rect 9518 22031 9590 22065
rect 9473 22021 9590 22031
rect 9245 21997 9590 22021
rect 9258 21953 9458 21997
rect 9473 21987 9497 21997
rect 9473 21963 9507 21987
rect 9518 21963 9590 21997
rect 9473 21953 9590 21963
rect 9245 21929 9590 21953
rect 9258 21885 9458 21929
rect 9473 21919 9497 21929
rect 9473 21895 9507 21919
rect 9518 21895 9590 21929
rect 9473 21885 9590 21895
rect 9245 21861 9590 21885
rect 9258 21817 9458 21861
rect 9473 21851 9497 21861
rect 9473 21827 9507 21851
rect 9518 21827 9590 21861
rect 9473 21817 9590 21827
rect 9245 21793 9590 21817
rect 9258 21749 9458 21793
rect 9473 21783 9497 21793
rect 9473 21759 9507 21783
rect 9518 21759 9590 21793
rect 9473 21749 9590 21759
rect 9245 21725 9590 21749
rect 9258 21681 9458 21725
rect 9473 21715 9497 21725
rect 9473 21691 9507 21715
rect 9518 21691 9590 21725
rect 9473 21681 9590 21691
rect 9245 21657 9590 21681
rect 9258 21613 9458 21657
rect 9473 21647 9497 21657
rect 9473 21623 9507 21647
rect 9518 21623 9590 21657
rect 9473 21613 9590 21623
rect 9245 21589 9590 21613
rect 9258 21545 9458 21589
rect 9473 21579 9497 21589
rect 9473 21555 9507 21579
rect 9518 21555 9590 21589
rect 9473 21545 9590 21555
rect 9245 21521 9590 21545
rect 9258 21477 9458 21521
rect 9473 21511 9497 21521
rect 9473 21487 9507 21511
rect 9518 21487 9590 21521
rect 9473 21477 9590 21487
rect 9245 21453 9590 21477
rect 9258 21409 9458 21453
rect 9473 21443 9497 21453
rect 9473 21419 9507 21443
rect 9518 21419 9590 21453
rect 9473 21409 9590 21419
rect 9245 21385 9590 21409
rect 9258 21315 9458 21385
rect 9473 21361 9497 21385
rect 9518 21315 9590 21385
rect 9820 21315 9876 22315
rect 9892 21315 9948 22315
rect 10250 22293 10450 22315
rect 10465 22303 10499 22327
rect 11253 22315 11287 22327
rect 10510 22303 10582 22315
rect 10465 22293 10582 22303
rect 10237 22269 10582 22293
rect 10250 22225 10450 22269
rect 10465 22259 10489 22269
rect 10465 22235 10499 22259
rect 10510 22235 10582 22269
rect 10465 22225 10582 22235
rect 10237 22201 10582 22225
rect 10250 22157 10450 22201
rect 10465 22191 10489 22201
rect 10465 22167 10499 22191
rect 10510 22167 10582 22201
rect 10465 22157 10582 22167
rect 10237 22133 10582 22157
rect 10250 22089 10450 22133
rect 10465 22123 10489 22133
rect 10465 22099 10499 22123
rect 10510 22099 10582 22133
rect 10465 22089 10582 22099
rect 10237 22065 10582 22089
rect 10250 22021 10450 22065
rect 10465 22055 10489 22065
rect 10465 22031 10499 22055
rect 10510 22031 10582 22065
rect 10465 22021 10582 22031
rect 10237 21997 10582 22021
rect 10250 21953 10450 21997
rect 10465 21987 10489 21997
rect 10465 21963 10499 21987
rect 10510 21963 10582 21997
rect 10465 21953 10582 21963
rect 10237 21929 10582 21953
rect 10250 21885 10450 21929
rect 10465 21919 10489 21929
rect 10465 21895 10499 21919
rect 10510 21895 10582 21929
rect 10465 21885 10582 21895
rect 10237 21861 10582 21885
rect 10250 21817 10450 21861
rect 10465 21851 10489 21861
rect 10465 21827 10499 21851
rect 10510 21827 10582 21861
rect 10465 21817 10582 21827
rect 10237 21793 10582 21817
rect 10250 21749 10450 21793
rect 10465 21783 10489 21793
rect 10465 21759 10499 21783
rect 10510 21759 10582 21793
rect 10465 21749 10582 21759
rect 10237 21725 10582 21749
rect 10250 21681 10450 21725
rect 10465 21715 10489 21725
rect 10465 21691 10499 21715
rect 10510 21691 10582 21725
rect 10465 21681 10582 21691
rect 10237 21657 10582 21681
rect 10250 21613 10450 21657
rect 10465 21647 10489 21657
rect 10465 21623 10499 21647
rect 10510 21623 10582 21657
rect 10465 21613 10582 21623
rect 10237 21589 10582 21613
rect 10250 21545 10450 21589
rect 10465 21579 10489 21589
rect 10465 21555 10499 21579
rect 10510 21555 10582 21589
rect 10465 21545 10582 21555
rect 10237 21521 10582 21545
rect 10250 21477 10450 21521
rect 10465 21511 10489 21521
rect 10465 21487 10499 21511
rect 10510 21487 10582 21521
rect 10465 21477 10582 21487
rect 10237 21453 10582 21477
rect 10250 21409 10450 21453
rect 10465 21443 10489 21453
rect 10465 21419 10499 21443
rect 10510 21419 10582 21453
rect 10465 21409 10582 21419
rect 10237 21385 10582 21409
rect 10250 21315 10450 21385
rect 10465 21361 10489 21385
rect 10510 21315 10582 21385
rect 10812 21315 10868 22315
rect 10884 21315 10940 22315
rect 11242 22293 11442 22315
rect 11457 22303 11491 22327
rect 12245 22315 12279 22327
rect 11502 22303 11574 22315
rect 11457 22293 11574 22303
rect 11229 22269 11574 22293
rect 11242 22225 11442 22269
rect 11457 22259 11481 22269
rect 11457 22235 11491 22259
rect 11502 22235 11574 22269
rect 11457 22225 11574 22235
rect 11229 22201 11574 22225
rect 11242 22157 11442 22201
rect 11457 22191 11481 22201
rect 11457 22167 11491 22191
rect 11502 22167 11574 22201
rect 11457 22157 11574 22167
rect 11229 22133 11574 22157
rect 11242 22089 11442 22133
rect 11457 22123 11481 22133
rect 11457 22099 11491 22123
rect 11502 22099 11574 22133
rect 11457 22089 11574 22099
rect 11229 22065 11574 22089
rect 11242 22021 11442 22065
rect 11457 22055 11481 22065
rect 11457 22031 11491 22055
rect 11502 22031 11574 22065
rect 11457 22021 11574 22031
rect 11229 21997 11574 22021
rect 11242 21953 11442 21997
rect 11457 21987 11481 21997
rect 11457 21963 11491 21987
rect 11502 21963 11574 21997
rect 11457 21953 11574 21963
rect 11229 21929 11574 21953
rect 11242 21885 11442 21929
rect 11457 21919 11481 21929
rect 11457 21895 11491 21919
rect 11502 21895 11574 21929
rect 11457 21885 11574 21895
rect 11229 21861 11574 21885
rect 11242 21817 11442 21861
rect 11457 21851 11481 21861
rect 11457 21827 11491 21851
rect 11502 21827 11574 21861
rect 11457 21817 11574 21827
rect 11229 21793 11574 21817
rect 11242 21749 11442 21793
rect 11457 21783 11481 21793
rect 11457 21759 11491 21783
rect 11502 21759 11574 21793
rect 11457 21749 11574 21759
rect 11229 21725 11574 21749
rect 11242 21681 11442 21725
rect 11457 21715 11481 21725
rect 11457 21691 11491 21715
rect 11502 21691 11574 21725
rect 11457 21681 11574 21691
rect 11229 21657 11574 21681
rect 11242 21613 11442 21657
rect 11457 21647 11481 21657
rect 11457 21623 11491 21647
rect 11502 21623 11574 21657
rect 11457 21613 11574 21623
rect 11229 21589 11574 21613
rect 11242 21545 11442 21589
rect 11457 21579 11481 21589
rect 11457 21555 11491 21579
rect 11502 21555 11574 21589
rect 11457 21545 11574 21555
rect 11229 21521 11574 21545
rect 11242 21477 11442 21521
rect 11457 21511 11481 21521
rect 11457 21487 11491 21511
rect 11502 21487 11574 21521
rect 11457 21477 11574 21487
rect 11229 21453 11574 21477
rect 11242 21409 11442 21453
rect 11457 21443 11481 21453
rect 11457 21419 11491 21443
rect 11502 21419 11574 21453
rect 11457 21409 11574 21419
rect 11229 21385 11574 21409
rect 11242 21315 11442 21385
rect 11457 21361 11481 21385
rect 11502 21315 11574 21385
rect 11804 21315 11860 22315
rect 11876 21315 11932 22315
rect 12234 22293 12434 22315
rect 12449 22303 12483 22327
rect 13237 22315 13271 22327
rect 12494 22303 12566 22315
rect 12449 22293 12566 22303
rect 12221 22269 12566 22293
rect 12234 22225 12434 22269
rect 12449 22259 12473 22269
rect 12449 22235 12483 22259
rect 12494 22235 12566 22269
rect 12449 22225 12566 22235
rect 12221 22201 12566 22225
rect 12234 22157 12434 22201
rect 12449 22191 12473 22201
rect 12449 22167 12483 22191
rect 12494 22167 12566 22201
rect 12449 22157 12566 22167
rect 12221 22133 12566 22157
rect 12234 22089 12434 22133
rect 12449 22123 12473 22133
rect 12449 22099 12483 22123
rect 12494 22099 12566 22133
rect 12449 22089 12566 22099
rect 12221 22065 12566 22089
rect 12234 22021 12434 22065
rect 12449 22055 12473 22065
rect 12449 22031 12483 22055
rect 12494 22031 12566 22065
rect 12449 22021 12566 22031
rect 12221 21997 12566 22021
rect 12234 21953 12434 21997
rect 12449 21987 12473 21997
rect 12449 21963 12483 21987
rect 12494 21963 12566 21997
rect 12449 21953 12566 21963
rect 12221 21929 12566 21953
rect 12234 21885 12434 21929
rect 12449 21919 12473 21929
rect 12449 21895 12483 21919
rect 12494 21895 12566 21929
rect 12449 21885 12566 21895
rect 12221 21861 12566 21885
rect 12234 21817 12434 21861
rect 12449 21851 12473 21861
rect 12449 21827 12483 21851
rect 12494 21827 12566 21861
rect 12449 21817 12566 21827
rect 12221 21793 12566 21817
rect 12234 21749 12434 21793
rect 12449 21783 12473 21793
rect 12449 21759 12483 21783
rect 12494 21759 12566 21793
rect 12449 21749 12566 21759
rect 12221 21725 12566 21749
rect 12234 21681 12434 21725
rect 12449 21715 12473 21725
rect 12449 21691 12483 21715
rect 12494 21691 12566 21725
rect 12449 21681 12566 21691
rect 12221 21657 12566 21681
rect 12234 21613 12434 21657
rect 12449 21647 12473 21657
rect 12449 21623 12483 21647
rect 12494 21623 12566 21657
rect 12449 21613 12566 21623
rect 12221 21589 12566 21613
rect 12234 21545 12434 21589
rect 12449 21579 12473 21589
rect 12449 21555 12483 21579
rect 12494 21555 12566 21589
rect 12449 21545 12566 21555
rect 12221 21521 12566 21545
rect 12234 21477 12434 21521
rect 12449 21511 12473 21521
rect 12449 21487 12483 21511
rect 12494 21487 12566 21521
rect 12449 21477 12566 21487
rect 12221 21453 12566 21477
rect 12234 21409 12434 21453
rect 12449 21443 12473 21453
rect 12449 21419 12483 21443
rect 12494 21419 12566 21453
rect 12449 21409 12566 21419
rect 12221 21385 12566 21409
rect 12234 21315 12434 21385
rect 12449 21361 12473 21385
rect 12494 21315 12566 21385
rect 12796 21315 12852 22315
rect 12868 21315 12924 22315
rect 13226 22293 13426 22315
rect 13441 22303 13475 22327
rect 14229 22315 14263 22327
rect 13486 22303 13558 22315
rect 13441 22293 13558 22303
rect 13213 22269 13558 22293
rect 13226 22225 13426 22269
rect 13441 22259 13465 22269
rect 13441 22235 13475 22259
rect 13486 22235 13558 22269
rect 13441 22225 13558 22235
rect 13213 22201 13558 22225
rect 13226 22157 13426 22201
rect 13441 22191 13465 22201
rect 13441 22167 13475 22191
rect 13486 22167 13558 22201
rect 13441 22157 13558 22167
rect 13213 22133 13558 22157
rect 13226 22089 13426 22133
rect 13441 22123 13465 22133
rect 13441 22099 13475 22123
rect 13486 22099 13558 22133
rect 13441 22089 13558 22099
rect 13213 22065 13558 22089
rect 13226 22021 13426 22065
rect 13441 22055 13465 22065
rect 13441 22031 13475 22055
rect 13486 22031 13558 22065
rect 13441 22021 13558 22031
rect 13213 21997 13558 22021
rect 13226 21953 13426 21997
rect 13441 21987 13465 21997
rect 13441 21963 13475 21987
rect 13486 21963 13558 21997
rect 13441 21953 13558 21963
rect 13213 21929 13558 21953
rect 13226 21885 13426 21929
rect 13441 21919 13465 21929
rect 13441 21895 13475 21919
rect 13486 21895 13558 21929
rect 13441 21885 13558 21895
rect 13213 21861 13558 21885
rect 13226 21817 13426 21861
rect 13441 21851 13465 21861
rect 13441 21827 13475 21851
rect 13486 21827 13558 21861
rect 13441 21817 13558 21827
rect 13213 21793 13558 21817
rect 13226 21749 13426 21793
rect 13441 21783 13465 21793
rect 13441 21759 13475 21783
rect 13486 21759 13558 21793
rect 13441 21749 13558 21759
rect 13213 21725 13558 21749
rect 13226 21681 13426 21725
rect 13441 21715 13465 21725
rect 13441 21691 13475 21715
rect 13486 21691 13558 21725
rect 13441 21681 13558 21691
rect 13213 21657 13558 21681
rect 13226 21613 13426 21657
rect 13441 21647 13465 21657
rect 13441 21623 13475 21647
rect 13486 21623 13558 21657
rect 13441 21613 13558 21623
rect 13213 21589 13558 21613
rect 13226 21545 13426 21589
rect 13441 21579 13465 21589
rect 13441 21555 13475 21579
rect 13486 21555 13558 21589
rect 13441 21545 13558 21555
rect 13213 21521 13558 21545
rect 13226 21477 13426 21521
rect 13441 21511 13465 21521
rect 13441 21487 13475 21511
rect 13486 21487 13558 21521
rect 13441 21477 13558 21487
rect 13213 21453 13558 21477
rect 13226 21409 13426 21453
rect 13441 21443 13465 21453
rect 13441 21419 13475 21443
rect 13486 21419 13558 21453
rect 13441 21409 13558 21419
rect 13213 21385 13558 21409
rect 13226 21315 13426 21385
rect 13441 21361 13465 21385
rect 13486 21315 13558 21385
rect 13788 21315 13844 22315
rect 13860 21315 13916 22315
rect 14218 22293 14418 22315
rect 14433 22303 14467 22327
rect 14478 22303 14550 22315
rect 14433 22293 14550 22303
rect 14205 22269 14550 22293
rect 14218 22225 14418 22269
rect 14433 22259 14457 22269
rect 14433 22235 14467 22259
rect 14478 22235 14550 22269
rect 14433 22225 14550 22235
rect 14205 22201 14550 22225
rect 14218 22157 14418 22201
rect 14433 22191 14457 22201
rect 14433 22167 14467 22191
rect 14478 22167 14550 22201
rect 14433 22157 14550 22167
rect 14205 22133 14550 22157
rect 14218 22089 14418 22133
rect 14433 22123 14457 22133
rect 14433 22099 14467 22123
rect 14478 22099 14550 22133
rect 14433 22089 14550 22099
rect 14205 22065 14550 22089
rect 14218 22021 14418 22065
rect 14433 22055 14457 22065
rect 14433 22031 14467 22055
rect 14478 22031 14550 22065
rect 14433 22021 14550 22031
rect 14205 21997 14550 22021
rect 14218 21953 14418 21997
rect 14433 21987 14457 21997
rect 14433 21963 14467 21987
rect 14478 21963 14550 21997
rect 14433 21953 14550 21963
rect 14205 21929 14550 21953
rect 14218 21885 14418 21929
rect 14433 21919 14457 21929
rect 14433 21895 14467 21919
rect 14478 21895 14550 21929
rect 14433 21885 14550 21895
rect 14205 21861 14550 21885
rect 14218 21817 14418 21861
rect 14433 21851 14457 21861
rect 14433 21827 14467 21851
rect 14478 21827 14550 21861
rect 14433 21817 14550 21827
rect 14205 21793 14550 21817
rect 14218 21749 14418 21793
rect 14433 21783 14457 21793
rect 14433 21759 14467 21783
rect 14478 21759 14550 21793
rect 14433 21749 14550 21759
rect 14205 21725 14550 21749
rect 14218 21681 14418 21725
rect 14433 21715 14457 21725
rect 14433 21691 14467 21715
rect 14478 21691 14550 21725
rect 14433 21681 14550 21691
rect 14205 21657 14550 21681
rect 14218 21613 14418 21657
rect 14433 21647 14457 21657
rect 14433 21623 14467 21647
rect 14478 21623 14550 21657
rect 14433 21613 14550 21623
rect 14205 21589 14550 21613
rect 14218 21545 14418 21589
rect 14433 21579 14457 21589
rect 14433 21555 14467 21579
rect 14478 21555 14550 21589
rect 14433 21545 14550 21555
rect 14205 21521 14550 21545
rect 14218 21477 14418 21521
rect 14433 21511 14457 21521
rect 14433 21487 14467 21511
rect 14478 21487 14550 21521
rect 14433 21477 14550 21487
rect 14205 21453 14550 21477
rect 14218 21409 14418 21453
rect 14433 21443 14457 21453
rect 14433 21419 14467 21443
rect 14478 21419 14550 21453
rect 14433 21409 14550 21419
rect 14205 21385 14550 21409
rect 14218 21315 14418 21385
rect 14433 21361 14457 21385
rect 14478 21315 14550 21385
rect 14739 21315 14811 22315
rect 14877 21315 14894 22315
rect 15064 21315 15097 22315
rect 828 20113 983 20203
rect 828 20077 7969 20113
rect 947 20046 983 20077
rect 1062 20046 1096 20070
rect 1130 20046 1164 20070
rect 1198 20046 1232 20070
rect 1266 20046 1300 20070
rect 1334 20046 1368 20070
rect 1402 20046 1436 20070
rect 1470 20046 1504 20070
rect 1538 20046 1572 20070
rect 1606 20046 1640 20070
rect 1674 20046 1708 20070
rect 1742 20046 1776 20070
rect 1810 20046 1844 20070
rect 1878 20046 1912 20070
rect 1946 20046 1980 20070
rect 2014 20046 2048 20070
rect 2082 20046 2116 20070
rect 2150 20046 2184 20070
rect 2218 20046 2252 20070
rect 2286 20046 2320 20070
rect 2354 20046 2388 20070
rect 2422 20046 2456 20070
rect 2490 20046 2524 20070
rect 2558 20046 2592 20070
rect 2626 20046 2660 20070
rect 2694 20046 2728 20070
rect 2762 20046 2796 20070
rect 2830 20046 2864 20070
rect 2898 20046 2932 20070
rect 2966 20046 3000 20070
rect 3034 20046 3068 20070
rect 3102 20046 3136 20070
rect 3170 20046 3204 20070
rect 3238 20046 3272 20070
rect 3306 20046 3340 20070
rect 3374 20046 3408 20070
rect 3442 20046 3476 20070
rect 3510 20046 3544 20070
rect 3578 20046 3612 20070
rect 3646 20046 3680 20070
rect 3714 20046 3748 20070
rect 3782 20046 3816 20070
rect 3850 20046 3884 20070
rect 3918 20046 3952 20070
rect 3986 20046 4020 20070
rect 4054 20046 4088 20070
rect 4122 20046 4156 20070
rect 4190 20046 4224 20070
rect 4258 20046 4292 20070
rect 4326 20046 4360 20070
rect 4394 20046 4428 20070
rect 4492 20046 4526 20070
rect 4560 20046 4594 20070
rect 4628 20046 4662 20070
rect 4696 20046 4730 20070
rect 4764 20046 4798 20070
rect 4832 20046 4866 20070
rect 4900 20046 4934 20070
rect 4968 20046 5002 20070
rect 5036 20046 5070 20070
rect 5104 20046 5138 20070
rect 5172 20046 5206 20070
rect 5240 20046 5274 20070
rect 5308 20046 5342 20070
rect 5376 20046 5410 20070
rect 5444 20046 5478 20070
rect 5512 20046 5546 20070
rect 5580 20046 5614 20070
rect 5648 20046 5682 20070
rect 5716 20046 5750 20070
rect 5784 20046 5818 20070
rect 5852 20046 5886 20070
rect 5920 20046 5954 20070
rect 5988 20046 6022 20070
rect 6056 20046 6090 20070
rect 6124 20046 6158 20070
rect 6192 20046 6226 20070
rect 6260 20046 6294 20070
rect 6328 20046 6362 20070
rect 6396 20046 6430 20070
rect 6464 20046 6498 20070
rect 6532 20046 6566 20070
rect 6600 20046 6634 20070
rect 6668 20046 6702 20070
rect 6736 20046 6770 20070
rect 6804 20046 6838 20070
rect 6872 20046 6906 20070
rect 6940 20046 6974 20070
rect 7008 20046 7042 20070
rect 7076 20046 7110 20070
rect 7144 20046 7178 20070
rect 7212 20046 7246 20070
rect 7280 20046 7314 20070
rect 7348 20046 7382 20070
rect 7416 20046 7450 20070
rect 7484 20046 7518 20070
rect 7552 20046 7586 20070
rect 7620 20046 7654 20070
rect 7688 20046 7722 20070
rect 7756 20046 7790 20070
rect 7824 20046 7858 20070
rect 7933 20046 7969 20077
rect 947 20023 7969 20046
rect 947 20010 1062 20023
rect 1096 20010 1130 20023
rect 1164 20010 1198 20023
rect 1232 20010 1266 20023
rect 1300 20010 1334 20023
rect 1368 20010 1402 20023
rect 1436 20010 1470 20023
rect 1504 20010 1538 20023
rect 1572 20010 1606 20023
rect 1640 20010 1674 20023
rect 1708 20010 1742 20023
rect 1776 20010 1810 20023
rect 1844 20010 1878 20023
rect 1912 20010 1946 20023
rect 1980 20010 2014 20023
rect 2048 20010 2082 20023
rect 2116 20010 2150 20023
rect 2184 20010 2218 20023
rect 2252 20010 2286 20023
rect 2320 20010 2354 20023
rect 2388 20010 2422 20023
rect 2456 20010 2490 20023
rect 2524 20010 2558 20023
rect 2592 20010 2626 20023
rect 2660 20010 2694 20023
rect 2728 20010 2762 20023
rect 2796 20010 2830 20023
rect 2864 20010 2898 20023
rect 2932 20010 2966 20023
rect 3000 20010 3034 20023
rect 3068 20010 3102 20023
rect 3136 20010 3170 20023
rect 3204 20010 3238 20023
rect 3272 20010 3306 20023
rect 3340 20010 3374 20023
rect 3408 20010 3442 20023
rect 3476 20010 3510 20023
rect 3544 20010 3578 20023
rect 3612 20010 3646 20023
rect 3680 20010 3714 20023
rect 3748 20010 3782 20023
rect 3816 20010 3850 20023
rect 3884 20010 3918 20023
rect 3952 20010 3986 20023
rect 4020 20010 4054 20023
rect 4088 20010 4122 20023
rect 4156 20010 4190 20023
rect 4224 20010 4258 20023
rect 4292 20010 4326 20023
rect 4360 20010 4394 20023
rect 4428 20010 4492 20023
rect 4526 20010 4560 20023
rect 4594 20010 4628 20023
rect 4662 20010 4696 20023
rect 4730 20010 4764 20023
rect 4798 20010 4832 20023
rect 4866 20010 4900 20023
rect 4934 20010 4968 20023
rect 5002 20010 5036 20023
rect 5070 20010 5104 20023
rect 5138 20010 5172 20023
rect 5206 20010 5240 20023
rect 5274 20010 5308 20023
rect 5342 20010 5376 20023
rect 5410 20010 5444 20023
rect 5478 20010 5512 20023
rect 5546 20010 5580 20023
rect 5614 20010 5648 20023
rect 5682 20010 5716 20023
rect 5750 20010 5784 20023
rect 5818 20010 5852 20023
rect 5886 20010 5920 20023
rect 5954 20010 5988 20023
rect 6022 20010 6056 20023
rect 6090 20010 6124 20023
rect 6158 20010 6192 20023
rect 6226 20010 6260 20023
rect 6294 20010 6328 20023
rect 6362 20010 6396 20023
rect 6430 20010 6464 20023
rect 6498 20010 6532 20023
rect 6566 20010 6600 20023
rect 6634 20010 6668 20023
rect 6702 20010 6736 20023
rect 6770 20010 6804 20023
rect 6838 20010 6872 20023
rect 6906 20010 6940 20023
rect 6974 20010 7008 20023
rect 7042 20010 7076 20023
rect 7110 20010 7144 20023
rect 7178 20010 7212 20023
rect 7246 20010 7280 20023
rect 7314 20010 7348 20023
rect 7382 20010 7416 20023
rect 7450 20010 7484 20023
rect 7518 20010 7552 20023
rect 7586 20010 7620 20023
rect 7654 20010 7688 20023
rect 7722 20010 7756 20023
rect 7790 20010 7824 20023
rect 7858 20010 7969 20023
rect 1749 19699 2749 19749
rect 2879 19699 4279 19749
rect 4641 19699 6041 19749
rect 6171 19699 7571 19749
rect 1749 19543 2749 19671
rect 2879 19543 4279 19671
rect 4641 19543 6041 19671
rect 6171 19543 7571 19671
rect 1749 19387 2749 19515
rect 2879 19387 4279 19515
rect 4641 19387 6041 19515
rect 6171 19387 7571 19515
rect 1749 19231 2749 19359
rect 2879 19231 4279 19359
rect 4641 19231 6041 19359
rect 6171 19231 7571 19359
rect 9582 19307 9752 19613
rect 12870 19277 12886 19343
rect 14894 19277 14910 19343
rect 1749 19081 2749 19131
rect 2879 19081 4279 19131
rect 4641 19081 6041 19131
rect 6171 19081 7571 19131
rect 1907 18644 1941 18668
rect 1975 18644 2009 18668
rect 2043 18644 2077 18668
rect 2111 18644 2145 18668
rect 2179 18644 2213 18668
rect 2247 18644 2281 18668
rect 2315 18644 2349 18668
rect 2383 18644 2417 18668
rect 2451 18644 2485 18668
rect 2519 18644 2553 18668
rect 2587 18644 2621 18668
rect 2655 18644 2689 18668
rect 2723 18644 2757 18668
rect 2791 18644 2825 18668
rect 2859 18644 2893 18668
rect 2927 18644 2961 18668
rect 2995 18644 3029 18668
rect 3063 18644 3097 18668
rect 3131 18644 3165 18668
rect 3199 18644 3233 18668
rect 3267 18644 3301 18668
rect 3335 18644 3369 18668
rect 3403 18644 3437 18668
rect 3471 18644 3505 18668
rect 3539 18644 3573 18668
rect 3607 18644 3641 18668
rect 3675 18644 3709 18668
rect 3743 18644 3777 18668
rect 3811 18644 3845 18668
rect 3879 18644 3913 18668
rect 3947 18644 3981 18668
rect 4015 18644 4049 18668
rect 4083 18644 4117 18668
rect 4151 18644 4185 18668
rect 4219 18644 4253 18668
rect 4287 18644 4321 18668
rect 4355 18644 4389 18668
rect 4423 18644 4457 18668
rect 4491 18644 4525 18668
rect 4559 18644 4593 18668
rect 4627 18644 4661 18668
rect 4695 18644 4729 18668
rect 4763 18644 4797 18668
rect 4831 18644 4865 18668
rect 4899 18644 4933 18668
rect 4967 18644 5001 18668
rect 5035 18644 5069 18668
rect 5103 18644 5137 18668
rect 5171 18644 5205 18668
rect 5239 18644 5273 18668
rect 5307 18644 5341 18668
rect 5375 18644 5409 18668
rect 5443 18644 5477 18668
rect 5511 18644 5545 18668
rect 5579 18644 5613 18668
rect 5647 18644 5681 18668
rect 5715 18653 5749 18668
rect 5697 18644 5749 18653
rect 5697 18619 5715 18644
rect 5731 18619 5749 18644
rect 5772 18619 5773 18644
rect 5731 18610 5773 18619
rect 2282 18280 5282 18330
rect 2282 18124 5282 18252
rect 5731 18208 5833 18232
rect 5731 18184 5755 18208
rect 5809 18184 5833 18208
rect 7214 18184 7248 18242
rect 7403 18208 7437 18242
rect 7475 18208 7509 18242
rect 7547 18208 7581 18242
rect 7619 18208 7653 18242
rect 7403 18184 7427 18208
rect 7629 18184 7653 18208
rect 7807 18208 7909 18232
rect 9037 18221 9061 18245
rect 8935 18208 8959 18211
rect 7807 18184 7831 18208
rect 7885 18184 7909 18208
rect 9013 18197 9037 18211
rect 9190 18208 9292 18232
rect 2282 17968 5282 18096
rect 2282 17812 5282 17940
rect 2282 17656 5282 17784
rect 2282 17500 5282 17628
rect 2282 17344 5282 17472
rect 2282 17194 5282 17244
rect 6119 16780 6162 18180
rect 6269 16780 6397 18180
rect 6432 16780 6560 18180
rect 6595 16780 6723 18180
rect 6758 16780 6886 18180
rect 6921 16780 7049 18180
rect 7084 16780 7127 18180
rect 7996 16780 8046 18180
rect 8153 16780 8281 18180
rect 8316 16780 8444 18180
rect 8479 16780 8607 18180
rect 8642 16780 8770 18180
rect 8805 16780 8848 18180
rect 8911 18163 8935 18187
rect 9037 18163 9061 18187
rect 9190 18184 9214 18208
rect 9268 18184 9292 18208
rect 2775 16381 2945 16687
rect 3575 16381 3745 16687
rect 4375 16381 4545 16687
rect 2775 15881 2945 16187
rect 3575 15881 3745 16187
rect 4375 15881 4545 16187
rect 232 14421 282 15021
rect 382 14421 510 15021
rect 538 14421 666 15021
rect 694 14421 750 15021
rect 850 14421 978 15021
rect 1006 14421 1134 15021
rect 1162 14421 1212 15021
rect 1292 14421 1342 15021
rect 1442 14421 1492 15021
rect 1930 14420 1980 15020
rect 2080 14420 2208 15020
rect 2236 14420 2364 15020
rect 2392 14420 2448 15020
rect 2548 14420 2676 15020
rect 2704 14420 2832 15020
rect 2860 14420 2910 15020
rect 2990 14420 3040 15020
rect 3140 14420 3190 15020
rect 3312 14420 3362 15020
rect 3462 14420 3512 15020
rect 3592 14420 3642 15020
rect 3742 14420 3870 15020
rect 3898 14420 4026 15020
rect 4054 14420 4110 15020
rect 4210 14420 4338 15020
rect 4366 14420 4494 15020
rect 4522 14420 4572 15020
rect 6119 14508 6162 15908
rect 6269 14508 6397 15908
rect 6432 14508 6560 15908
rect 6595 14508 6723 15908
rect 6758 14508 6886 15908
rect 6921 14508 7049 15908
rect 7084 14508 7127 15908
rect 5731 14480 5833 14504
rect 5809 14456 5833 14480
rect 7214 14456 7248 14514
rect 7403 14480 7437 14514
rect 7475 14480 7509 14514
rect 7547 14480 7581 14514
rect 7619 14480 7653 14514
rect 7996 14508 8046 15908
rect 8153 14508 8281 15908
rect 8316 14508 8444 15908
rect 8479 14508 8607 15908
rect 8642 14508 8770 15908
rect 8805 14508 8848 15908
rect 7403 14456 7427 14480
rect 7629 14456 7653 14480
rect 7807 14480 7909 14504
rect 8911 14501 8935 14525
rect 9037 14501 9061 14525
rect 7807 14456 7831 14480
rect 7885 14456 7909 14480
rect 8935 14477 8959 14480
rect 9013 14477 9037 14491
rect 9190 14480 9292 14504
rect 9037 14443 9061 14467
rect 9190 14456 9214 14480
rect 9268 14456 9292 14480
rect 9468 14040 10004 18648
rect 12439 18340 12530 18442
rect 12763 18407 12777 18431
rect 12729 18383 12753 18407
rect 12787 18383 12811 18407
rect 15983 18333 16017 18353
rect 12386 18220 12410 18244
rect 12444 18220 12468 18244
rect 12920 18238 12954 18242
rect 12988 18238 13022 18242
rect 13056 18238 13090 18242
rect 13124 18238 13158 18242
rect 13192 18238 13226 18242
rect 13260 18238 13294 18242
rect 13328 18238 13362 18242
rect 13396 18238 13430 18242
rect 13464 18238 13498 18242
rect 13532 18238 13566 18242
rect 13600 18238 13634 18242
rect 13668 18238 13702 18242
rect 13736 18238 13770 18242
rect 13804 18238 13838 18242
rect 13872 18238 13906 18242
rect 13940 18238 13974 18242
rect 14008 18238 14042 18242
rect 14076 18238 14110 18242
rect 14144 18238 14178 18242
rect 14212 18238 14246 18242
rect 14280 18238 14314 18242
rect 14348 18238 14382 18242
rect 14416 18238 14450 18242
rect 14484 18238 14518 18242
rect 14552 18238 14586 18242
rect 14620 18238 14654 18242
rect 14688 18238 14722 18242
rect 14756 18238 14790 18242
rect 14824 18238 14858 18242
rect 14892 18238 14926 18242
rect 14960 18238 14994 18242
rect 15028 18238 15062 18242
rect 15096 18238 15130 18242
rect 15164 18238 15198 18242
rect 15232 18238 15266 18242
rect 15300 18238 15334 18242
rect 15368 18238 15402 18242
rect 15436 18238 15470 18242
rect 15504 18238 15538 18242
rect 15572 18238 15606 18242
rect 15640 18238 15674 18242
rect 12852 18220 15752 18238
rect 12920 18216 12954 18220
rect 12988 18216 13022 18220
rect 13056 18216 13090 18220
rect 13124 18216 13158 18220
rect 13192 18216 13226 18220
rect 13260 18216 13294 18220
rect 13328 18216 13362 18220
rect 13396 18216 13430 18220
rect 13464 18216 13498 18220
rect 13532 18216 13566 18220
rect 13600 18216 13634 18220
rect 13668 18216 13702 18220
rect 13736 18216 13770 18220
rect 13804 18216 13838 18220
rect 13872 18216 13906 18220
rect 13940 18216 13974 18220
rect 14008 18216 14042 18220
rect 14076 18216 14110 18220
rect 14144 18216 14178 18220
rect 14212 18216 14246 18220
rect 14280 18216 14314 18220
rect 14348 18216 14382 18220
rect 14416 18216 14450 18220
rect 14484 18216 14518 18220
rect 14552 18216 14586 18220
rect 14620 18216 14654 18220
rect 14688 18216 14722 18220
rect 14756 18216 14790 18220
rect 14824 18216 14858 18220
rect 14892 18216 14926 18220
rect 14960 18216 14994 18220
rect 15028 18216 15062 18220
rect 15096 18216 15130 18220
rect 15164 18216 15198 18220
rect 15232 18216 15266 18220
rect 15300 18216 15334 18220
rect 15368 18216 15402 18220
rect 15436 18216 15470 18220
rect 15504 18216 15538 18220
rect 15572 18216 15606 18220
rect 15640 18216 15674 18220
rect 15891 18217 15915 18241
rect 12410 18196 12444 18210
rect 12856 18208 15748 18216
rect 12896 18196 15698 18208
rect 15915 18193 15939 18208
rect 15983 18197 16017 18232
rect 10038 16780 10166 18180
rect 10201 16780 10329 18180
rect 10364 16780 10492 18180
rect 10527 16780 10655 18180
rect 10690 16780 10818 18180
rect 10853 16780 10981 18180
rect 11016 16780 11059 18180
rect 11152 16780 11195 18180
rect 11302 16780 11430 18180
rect 11465 16780 11593 18180
rect 11628 16780 11756 18180
rect 11791 16780 11919 18180
rect 11954 16780 12082 18180
rect 12117 16780 12245 18180
rect 12280 16780 12330 18180
rect 12386 18162 12410 18186
rect 12444 18162 12468 18186
rect 15993 18184 16017 18197
rect 12597 16395 12699 17959
rect 12966 16712 13016 18112
rect 13123 16712 13251 18112
rect 13286 16712 13414 18112
rect 13449 16712 13577 18112
rect 13612 16712 13740 18112
rect 13775 16712 13903 18112
rect 13938 16712 14066 18112
rect 14101 16712 14144 18112
rect 14237 16712 14280 18112
rect 14387 16712 14515 18112
rect 14550 16712 14678 18112
rect 14713 16712 14841 18112
rect 14876 16712 15004 18112
rect 15039 16712 15167 18112
rect 15202 16712 15330 18112
rect 15365 16712 15493 18112
rect 15528 16712 15571 18112
rect 12631 16371 12665 16395
rect 12631 16293 12665 16317
rect 10038 14508 10166 15908
rect 10201 14508 10329 15908
rect 10364 14508 10492 15908
rect 10527 14508 10655 15908
rect 10690 14508 10818 15908
rect 10853 14508 10981 15908
rect 11016 14508 11059 15908
rect 11152 14508 11195 15908
rect 11302 14508 11430 15908
rect 11465 14508 11593 15908
rect 11628 14508 11756 15908
rect 11791 14508 11919 15908
rect 11954 14508 12082 15908
rect 12117 14508 12245 15908
rect 12280 14508 12330 15908
rect 12597 14729 12699 16293
rect 12966 14576 13016 15976
rect 13123 14576 13251 15976
rect 13286 14576 13414 15976
rect 13449 14576 13577 15976
rect 13612 14576 13740 15976
rect 13775 14576 13903 15976
rect 13938 14576 14066 15976
rect 14101 14576 14144 15976
rect 14237 14576 14280 15976
rect 14387 14576 14515 15976
rect 14550 14576 14678 15976
rect 14713 14576 14841 15976
rect 14876 14576 15004 15976
rect 15039 14576 15167 15976
rect 15202 14576 15330 15976
rect 15365 14576 15493 15976
rect 15528 14576 15571 15976
rect 12386 14502 12410 14526
rect 12444 14502 12468 14526
rect 12920 14510 12954 14514
rect 12988 14510 13022 14514
rect 13056 14510 13090 14514
rect 13124 14510 13158 14514
rect 13192 14510 13226 14514
rect 13260 14510 13294 14514
rect 13328 14510 13362 14514
rect 13396 14510 13430 14514
rect 13464 14510 13498 14514
rect 13532 14510 13566 14514
rect 13600 14510 13634 14514
rect 13668 14510 13702 14514
rect 13736 14510 13770 14514
rect 13804 14510 13838 14514
rect 13872 14510 13906 14514
rect 13940 14510 13974 14514
rect 14008 14510 14042 14514
rect 14076 14510 14110 14514
rect 14144 14510 14178 14514
rect 14212 14510 14246 14514
rect 14280 14510 14314 14514
rect 14348 14510 14382 14514
rect 14416 14510 14450 14514
rect 14484 14510 14518 14514
rect 14552 14510 14586 14514
rect 14620 14510 14654 14514
rect 14688 14510 14722 14514
rect 14756 14510 14790 14514
rect 14824 14510 14858 14514
rect 14892 14510 14926 14514
rect 14960 14510 14994 14514
rect 15028 14510 15062 14514
rect 15096 14510 15130 14514
rect 15164 14510 15198 14514
rect 15232 14510 15266 14514
rect 15300 14510 15334 14514
rect 15368 14510 15402 14514
rect 15436 14510 15470 14514
rect 15504 14510 15538 14514
rect 15572 14510 15606 14514
rect 15640 14510 15674 14514
rect 12886 14502 15718 14510
rect 15949 14505 16017 14525
rect 12920 14498 12954 14502
rect 12988 14498 13022 14502
rect 13056 14498 13090 14502
rect 13124 14498 13158 14502
rect 13192 14498 13226 14502
rect 13260 14498 13294 14502
rect 13328 14498 13362 14502
rect 13396 14498 13430 14502
rect 13464 14498 13498 14502
rect 13532 14498 13566 14502
rect 13600 14498 13634 14502
rect 13668 14498 13702 14502
rect 13736 14498 13770 14502
rect 13804 14498 13838 14502
rect 13872 14498 13906 14502
rect 13940 14498 13974 14502
rect 14008 14498 14042 14502
rect 14076 14498 14110 14502
rect 14144 14498 14178 14502
rect 14212 14498 14246 14502
rect 14280 14498 14314 14502
rect 14348 14498 14382 14502
rect 14416 14498 14450 14502
rect 14484 14498 14518 14502
rect 14552 14498 14586 14502
rect 14620 14498 14654 14502
rect 14688 14498 14722 14502
rect 14756 14498 14790 14502
rect 14824 14498 14858 14502
rect 14892 14498 14926 14502
rect 14960 14498 14994 14502
rect 15028 14498 15062 14502
rect 15096 14498 15130 14502
rect 15164 14498 15198 14502
rect 15232 14498 15266 14502
rect 15300 14498 15334 14502
rect 15368 14498 15402 14502
rect 15436 14498 15470 14502
rect 15504 14498 15538 14502
rect 15572 14498 15606 14502
rect 15640 14498 15674 14502
rect 12410 14478 12444 14492
rect 12852 14480 15752 14498
rect 15915 14480 15939 14495
rect 15983 14480 16017 14505
rect 12896 14478 15698 14480
rect 12386 14444 12410 14468
rect 12444 14444 12468 14468
rect 15891 14447 15915 14471
rect 15993 14456 16017 14480
rect 15949 14369 16017 14389
rect 12439 14246 12530 14348
rect 12729 14281 12753 14305
rect 12787 14281 12811 14305
rect 12763 14257 12777 14281
rect 2628 12903 2678 13103
rect 2778 12903 2834 13103
rect 2934 12903 2984 13103
rect 3334 12903 3384 13103
rect 3484 12903 3540 13103
rect 3640 12903 3690 13103
rect 3754 12903 3765 13103
rect 10618 12657 10668 13657
rect 10768 12657 10824 13657
rect 10924 12657 10980 13657
rect 11080 12657 11136 13657
rect 11236 13200 11286 13657
rect 11700 13200 11750 13657
rect 11236 13116 11289 13200
rect 11697 13116 11750 13200
rect 11236 12867 11286 13116
rect 11700 12867 11750 13116
rect 11236 12783 11289 12867
rect 11697 12783 11750 12867
rect 11236 12657 11286 12783
rect 11700 12657 11750 12783
rect 11850 12657 11906 13657
rect 12006 12657 12062 13657
rect 12162 12657 12218 13657
rect 12318 12657 12368 13657
rect 14553 13268 14603 13868
rect 14703 13268 14753 13868
rect 14825 13268 14875 13868
rect 14975 13268 15025 13868
rect 15101 13268 15151 13868
rect 15251 13268 15301 13868
rect 15373 13268 15423 13868
rect 15523 13268 15573 13868
rect 13509 12945 13815 13115
rect 10767 12319 10817 12435
rect 10764 12235 10817 12319
rect 10937 12235 11065 12435
rect 11113 12235 11169 12435
rect 11289 12235 11417 12435
rect 11465 12235 11521 12435
rect 11641 12235 11769 12435
rect 11817 12235 11873 12435
rect 11993 12235 12121 12435
rect 12169 12319 12219 12435
rect 14630 12381 15630 12431
rect 12169 12235 12222 12319
rect 10772 12231 10806 12235
rect 12180 12231 12214 12235
rect 14630 12225 15630 12353
rect 14630 12069 15630 12197
rect 10705 11921 11705 11971
rect 12897 11921 13897 11971
rect 14630 11913 15630 12041
rect 3068 11302 3118 11902
rect 3218 11302 3268 11902
rect 3348 11302 3398 11902
rect 3498 11302 3626 11902
rect 3654 11302 3782 11902
rect 3810 11302 3866 11902
rect 3966 11302 4094 11902
rect 4122 11302 4250 11902
rect 4278 11302 4328 11902
rect 10705 11765 11705 11821
rect 12897 11765 13897 11821
rect 14630 11757 15630 11885
rect 12043 11681 12127 11684
rect 10705 11609 11705 11665
rect 11927 11631 12127 11681
rect 12475 11681 12559 11684
rect 12475 11676 12675 11681
rect 12471 11642 12675 11676
rect 12475 11631 12675 11642
rect 12897 11609 13897 11665
rect 14630 11601 15630 11729
rect 10705 11453 11705 11509
rect 11927 11455 12127 11583
rect 12475 11455 12675 11583
rect 12897 11453 13897 11509
rect 14630 11445 15630 11573
rect 10705 11297 11705 11353
rect 11927 11279 12127 11335
rect 12475 11279 12675 11335
rect 12897 11297 13897 11353
rect 14630 11289 15630 11417
rect 10705 11147 11705 11197
rect 11163 11144 11247 11147
rect 11495 11144 11579 11147
rect 11927 11103 12127 11231
rect 12475 11103 12675 11231
rect 12897 11147 13897 11197
rect 13023 11144 13107 11147
rect 13355 11144 13439 11147
rect 14630 11133 15630 11261
rect 6369 10910 6403 10944
rect 6438 10910 6472 10944
rect 6507 10910 6541 10944
rect 6576 10910 6610 10944
rect 6645 10910 6679 10944
rect 6714 10910 6748 10944
rect 6783 10910 6817 10944
rect 6852 10910 6886 10944
rect 6921 10910 6955 10944
rect 6990 10910 7024 10944
rect 7059 10910 7093 10944
rect 7128 10910 7162 10944
rect 7197 10910 7231 10944
rect 7266 10910 7300 10944
rect 7335 10910 7369 10944
rect 7404 10910 7438 10944
rect 7473 10910 7507 10944
rect 7542 10910 7576 10944
rect 7611 10910 7645 10944
rect 7680 10910 7714 10944
rect 7749 10910 7783 10944
rect 7818 10910 7852 10944
rect 7887 10910 7921 10944
rect 7956 10910 7990 10944
rect 8025 10910 8059 10944
rect 8094 10910 8128 10944
rect 8163 10910 8197 10944
rect 8232 10910 8266 10944
rect 8301 10910 8335 10944
rect 8370 10910 8404 10944
rect 8439 10911 8468 10944
rect 11927 10933 12127 10983
rect 12475 10933 12675 10983
rect 14630 10977 15630 11105
rect 8439 10910 8502 10911
rect 6369 10886 6393 10910
rect 14630 10821 15630 10949
rect 14630 10665 15630 10793
rect 14630 10509 15630 10637
rect 14630 10353 15630 10481
rect 14630 10203 15630 10253
rect 9081 9791 9105 9815
rect 9141 9791 9165 9815
rect 11456 9791 11480 9815
rect 11515 9791 11539 9815
rect 9117 9767 9129 9791
rect 11491 9767 11504 9791
rect 9119 9703 9153 9713
rect 9095 9679 9153 9703
rect 11501 9679 11535 9713
rect 12128 9703 12162 9713
rect 12104 9679 12162 9703
rect 13838 9678 13862 9702
rect 13767 9662 13838 9668
rect 13814 9654 13838 9662
rect 1955 8822 2005 9422
rect 2125 8822 2181 9422
rect 2301 8822 2351 9422
rect 656 8736 680 8760
rect 717 8750 741 8760
rect 717 8746 751 8750
rect 788 8746 822 8750
rect 859 8746 893 8750
rect 695 8736 917 8746
rect 693 8732 704 8736
rect 717 8732 751 8736
rect 788 8732 822 8736
rect 859 8732 893 8736
rect 693 8712 917 8732
rect 717 8692 741 8712
rect 2440 8600 2490 9600
rect 2590 8600 2640 9600
rect 2749 8600 2799 9600
rect 2899 8600 2949 9600
rect 3079 9140 3259 9340
rect 3424 9325 3484 9340
rect 3510 9325 3570 9340
rect 5084 9325 5144 9340
rect 5170 9325 5230 9340
rect 3439 9155 3469 9325
rect 3525 9155 3555 9325
rect 5099 9155 5129 9325
rect 5185 9155 5215 9325
rect 3428 9152 3480 9155
rect 3514 9152 3566 9155
rect 5088 9152 5140 9155
rect 5174 9152 5226 9155
rect 3424 9140 3484 9152
rect 3510 9140 3570 9152
rect 5084 9140 5144 9152
rect 5170 9140 5230 9152
rect 5395 9140 5575 9340
rect 3079 8880 3259 9080
rect 3424 9065 3484 9080
rect 3510 9065 3570 9080
rect 5084 9065 5144 9080
rect 5170 9065 5230 9080
rect 3439 8895 3469 9065
rect 3525 8895 3555 9065
rect 5099 8895 5129 9065
rect 5185 8895 5215 9065
rect 3428 8892 3480 8895
rect 3514 8892 3566 8895
rect 5088 8892 5140 8895
rect 5174 8892 5226 8895
rect 3424 8880 3484 8892
rect 3510 8880 3570 8892
rect 5084 8880 5144 8892
rect 5170 8880 5230 8892
rect 5395 8880 5575 9080
rect 3079 8620 3259 8820
rect 3424 8805 3484 8820
rect 3510 8805 3570 8820
rect 5084 8805 5144 8820
rect 5170 8805 5230 8820
rect 3439 8800 3469 8805
rect 3525 8800 3555 8805
rect 5099 8800 5129 8805
rect 5185 8800 5215 8805
rect 5395 8620 5575 8820
rect 5705 8600 5755 9600
rect 5855 8600 5905 9600
rect 6014 8600 6064 9600
rect 6164 8600 6214 9600
rect 7528 9566 13277 9578
rect 6303 8822 6353 9422
rect 6473 8822 6529 9422
rect 6649 8822 6699 9422
rect 7528 8875 7554 9566
rect 7544 8872 7554 8875
rect 7688 8858 7738 9458
rect 7858 8858 7914 9458
rect 8034 8858 8084 9458
rect 8150 8858 8200 9458
rect 8320 8858 8376 9458
rect 8496 8858 8624 9458
rect 8672 8858 8800 9458
rect 8848 8858 8976 9458
rect 9024 8858 9074 9458
rect 9140 8858 9190 9458
rect 9310 8858 9438 9458
rect 9486 8858 9542 9458
rect 9662 8858 9790 9458
rect 9838 8858 9888 9458
rect 9954 8858 10004 9458
rect 10124 8858 10252 9458
rect 10300 8858 10428 9458
rect 10476 8858 10604 9458
rect 10652 8858 10780 9458
rect 10828 8858 10956 9458
rect 11004 8858 11060 9458
rect 11180 8858 11308 9458
rect 11356 8858 11484 9458
rect 11532 8858 11660 9458
rect 11708 8858 11836 9458
rect 11884 8858 12012 9458
rect 12060 8858 12116 9458
rect 12236 8858 12364 9458
rect 12412 8858 12468 9458
rect 12588 8858 12716 9458
rect 12764 8858 12820 9458
rect 12940 8858 13068 9458
rect 13116 8858 13166 9458
rect 14591 9148 14771 9348
rect 14827 9148 15007 9348
rect 14591 9013 14771 9050
rect 15278 8748 15328 9348
rect 15448 8748 15504 9348
rect 15624 8748 15680 9348
rect 15800 8748 15850 9348
rect 3079 8306 3259 8506
rect 5395 8306 5575 8506
rect 1443 7530 1493 8130
rect 1593 7530 1649 8130
rect 1749 7530 1799 8130
rect 2483 8046 2663 8246
rect 2719 8046 2899 8246
rect 3079 8046 3259 8246
rect 3424 8231 3484 8246
rect 3510 8231 3570 8246
rect 5084 8231 5144 8246
rect 5170 8231 5230 8246
rect 3439 8061 3469 8231
rect 3525 8061 3555 8231
rect 3428 8058 3480 8061
rect 3514 8058 3566 8061
rect 3424 8046 3484 8058
rect 3510 8046 3570 8058
rect 2483 7786 2663 7986
rect 2719 7786 2899 7986
rect 3079 7786 3259 7986
rect 3424 7971 3484 7986
rect 3510 7971 3570 7986
rect 3439 7801 3469 7971
rect 3525 7801 3555 7971
rect 3428 7798 3480 7801
rect 3514 7798 3566 7801
rect 3424 7786 3484 7798
rect 3510 7786 3570 7798
rect 3716 7796 3732 8112
rect 4920 7796 4938 8112
rect 5099 8061 5129 8231
rect 5185 8061 5215 8231
rect 5088 8058 5140 8061
rect 5174 8058 5226 8061
rect 5084 8046 5144 8058
rect 5170 8046 5230 8058
rect 5395 8046 5575 8246
rect 5755 8046 5935 8246
rect 5991 8046 6171 8246
rect 5084 7971 5144 7986
rect 5170 7971 5230 7986
rect 5099 7801 5129 7971
rect 5185 7801 5215 7971
rect 5088 7798 5140 7801
rect 5174 7798 5226 7801
rect 3716 7770 3720 7796
rect 5084 7786 5144 7798
rect 5170 7786 5230 7798
rect 5395 7786 5575 7986
rect 5755 7786 5935 7986
rect 5991 7786 6171 7986
rect 3079 7526 3259 7726
rect 3424 7711 3484 7726
rect 3510 7711 3570 7726
rect 3439 7672 3469 7711
rect 3525 7672 3555 7711
rect 3682 7532 3720 7770
rect 4940 7532 4972 7770
rect 5084 7711 5144 7726
rect 5170 7711 5230 7726
rect 5099 7672 5129 7711
rect 5185 7672 5215 7711
rect 5395 7526 5575 7726
rect 6855 7530 6905 8130
rect 7005 7530 7061 8130
rect 7161 7530 7211 8130
rect 7708 7544 7758 8544
rect 7858 7544 7914 8544
rect 8014 7544 8064 8544
rect 8150 7544 8200 8544
rect 8300 7544 8356 8544
rect 8456 7544 8512 8544
rect 8612 7544 8668 8544
rect 8768 7544 8818 8544
rect 8884 7544 8934 8544
rect 9034 7544 9162 8544
rect 9190 7544 9318 8544
rect 9346 7544 9474 8544
rect 9502 7544 9630 8544
rect 9658 7544 9786 8544
rect 9814 7544 9870 8544
rect 9970 7544 10098 8544
rect 10126 7544 10254 8544
rect 10282 7544 10410 8544
rect 10438 7544 10566 8544
rect 10594 7544 10722 8544
rect 10750 7544 10806 8544
rect 10926 7544 11054 8544
rect 11102 7544 11230 8544
rect 11278 7544 11406 8544
rect 11454 7544 11582 8544
rect 11630 7544 11758 8544
rect 11806 7544 11934 8544
rect 11982 7544 12110 8544
rect 12158 7544 12208 8544
rect 12274 7544 12324 8544
rect 12424 7544 12552 8544
rect 12580 7544 12708 8544
rect 12736 7544 12864 8544
rect 12892 7544 12948 8544
rect 13048 7544 13176 8544
rect 13204 7544 13332 8544
rect 13360 7544 13488 8544
rect 13516 7544 13566 8544
rect 14157 7985 14210 8135
rect 14160 7888 14210 7985
rect 14157 7666 14210 7888
rect 14160 7535 14210 7666
rect 14330 7535 14386 8135
rect 14506 7535 14556 8135
rect 14932 7540 14982 8140
rect 15102 7540 15152 8140
rect 160 6558 168 6783
rect 237 5701 287 6301
rect 387 5701 437 6301
rect 1293 6063 1343 6663
rect 1443 6063 1499 6663
rect 1599 6063 1649 6663
rect 1821 5997 1871 6997
rect 1971 5997 2027 6997
rect 2127 5997 2177 6997
rect 2243 5997 2293 6997
rect 2393 5997 2521 6997
rect 2549 5997 2677 6997
rect 2705 5997 2833 6997
rect 2861 5997 2917 6997
rect 3017 5997 3145 6997
rect 3173 5997 3301 6997
rect 3329 5997 3457 6997
rect 3485 5997 3535 6997
rect 3687 5997 3737 6997
rect 3837 5997 3965 6997
rect 3993 5997 4121 6997
rect 4149 5997 4277 6997
rect 4305 5997 4433 6997
rect 4461 5997 4589 6997
rect 4617 5997 4745 6997
rect 4773 5997 4901 6997
rect 4929 5997 4979 6997
rect 5131 6047 5181 7047
rect 5281 6047 5409 7047
rect 5437 6047 5565 7047
rect 5593 6047 5721 7047
rect 5749 6047 5877 7047
rect 5905 6047 6033 7047
rect 6061 6047 6189 7047
rect 6217 6047 6345 7047
rect 6373 6047 6423 7047
rect 6575 5997 6625 6997
rect 6725 5997 6853 6997
rect 6881 5997 7009 6997
rect 7037 5997 7165 6997
rect 7193 5997 7321 6997
rect 7349 5997 7477 6997
rect 7505 5997 7633 6997
rect 7661 5997 7789 6997
rect 7817 5997 7873 6997
rect 7973 5997 8023 6997
rect 8175 6397 8225 6997
rect 8609 6397 8659 6997
rect 9852 6512 9902 7112
rect 10002 6512 10130 7112
rect 10158 6512 10286 7112
rect 10314 6512 10364 7112
rect 10444 6512 10494 7112
rect 10594 6512 10722 7112
rect 10750 6512 10806 7112
rect 10906 6512 11034 7112
rect 11062 6512 11112 7112
rect 11192 6512 11242 7112
rect 11342 6512 11398 7112
rect 11498 6512 11548 7112
rect 10477 5732 10513 6332
rect 10837 5732 10893 6332
rect 11027 5732 11077 6332
rect 6740 5618 6806 5634
rect 6902 5618 6968 5634
rect 9310 5564 9385 5574
rect 9605 5564 9680 5574
rect 1593 4914 1643 5514
rect 1743 4914 1799 5514
rect 1899 4914 1949 5514
rect 2161 4883 2211 5483
rect 2311 4883 2439 5483
rect 2467 4883 2595 5483
rect 2623 4883 2751 5483
rect 2779 4883 2829 5483
rect 2895 4883 2945 5483
rect 3045 4883 3173 5483
rect 3201 4883 3329 5483
rect 3357 4883 3485 5483
rect 3513 4883 3569 5483
rect 3669 4883 3797 5483
rect 3825 4883 3953 5483
rect 3981 4883 4109 5483
rect 4137 4883 4193 5483
rect 4293 4883 4349 5483
rect 4449 4883 4505 5483
rect 4605 4883 4655 5483
rect 4721 4883 4771 5483
rect 4871 4883 4999 5483
rect 5027 4883 5083 5483
rect 5183 4883 5311 5483
rect 5339 4883 5389 5483
rect 8322 5391 9322 5441
rect 9385 5391 9435 5502
rect 9382 5271 9435 5391
rect 8322 5221 9322 5271
rect 8285 4501 8335 5101
rect 8455 4501 8511 5101
rect 8631 4501 8681 5101
rect 8901 4502 8951 5102
rect 9071 4502 9127 5102
rect 9247 4502 9297 5102
rect 9385 4502 9435 5271
rect 9555 4502 9605 5502
rect 9668 5391 10268 5441
rect 9668 5291 9680 5391
rect 11567 5321 11617 5921
rect 11737 5321 11793 5921
rect 11913 5321 12041 5921
rect 12089 5321 12145 5921
rect 12265 5321 12321 5921
rect 12441 5321 12497 5921
rect 12617 5321 12745 5921
rect 12793 5321 12843 5921
rect 9668 5241 10268 5291
rect 9684 4502 9734 5102
rect 9854 4502 9910 5102
rect 10030 4502 10080 5102
rect 10371 4502 10421 5102
rect 10541 4502 10669 5102
rect 10717 4502 10773 5102
rect 10893 4502 11021 5102
rect 11069 4502 11119 5102
rect 11491 4566 11541 5166
rect 11661 4566 11789 5166
rect 11837 4566 11965 5166
rect 12013 4566 12141 5166
rect 12189 4566 12317 5166
rect 12365 4566 12421 5166
rect 12541 4566 12669 5166
rect 12717 4566 12767 5166
rect 4168 4378 4218 4459
rect 501 4047 516 4062
rect 465 4017 516 4047
rect 501 4002 516 4017
rect 1359 3706 1409 4306
rect 1529 3706 1657 4306
rect 1705 3706 1761 4306
rect 1881 3877 1931 4306
rect 1994 4106 2006 4306
rect 4165 4106 4218 4378
rect 1881 3805 1934 3877
rect 4168 3859 4218 4106
rect 4318 3859 4368 4459
rect 4434 3859 4484 4459
rect 4584 3859 4712 4459
rect 4740 3859 4868 4459
rect 4896 3859 5024 4459
rect 5102 3859 5155 4459
rect 1881 3706 1931 3805
rect 1994 3706 2006 3805
rect 4505 3495 4995 3522
rect 5105 3459 5155 3859
rect 5255 3459 5383 4459
rect 5411 3459 5461 4459
rect 5662 3338 5674 4338
rect 5731 3338 5781 4338
rect 5901 3338 6029 4338
rect 6077 3338 6205 4338
rect 6253 3338 6309 4338
rect 6429 3338 6479 4338
rect 6578 4218 6644 4234
rect 7064 4218 7130 4234
rect 6578 3434 6644 3450
rect 6740 3434 6806 3450
rect 6902 3434 6968 3450
rect 7064 3434 7130 3450
rect 7229 3338 7279 4338
rect 7399 3338 7455 4338
rect 7575 3338 7703 4338
rect 7751 3338 7879 4338
rect 7927 3338 7977 4338
rect 8034 3338 8046 4338
rect 8070 4274 8080 4308
rect 8070 4206 8080 4240
rect 8070 4138 8080 4172
rect 8070 4070 8080 4104
rect 8070 3995 8080 4029
rect 8070 3927 8080 3961
rect 8070 3859 8080 3893
rect 8070 3791 8080 3825
rect 8070 3723 8080 3757
rect 8070 3655 8080 3689
rect 8070 3587 8080 3621
rect 8070 3519 8080 3553
rect 8070 3451 8080 3485
rect 8070 3383 8080 3417
rect 8129 3338 8179 4338
rect 8299 3338 8427 4338
rect 8475 3338 8531 4338
rect 8651 3338 8701 4338
rect 8867 3738 8917 4338
rect 9037 3738 9093 4338
rect 9213 3738 9341 4338
rect 9389 3738 9439 4338
rect 9591 3738 9641 4338
rect 9741 3738 9869 4338
rect 9897 3738 9953 4338
rect 10053 3738 10181 4338
rect 10209 3738 10259 4338
rect 10463 3738 10513 4338
rect 10613 3738 10741 4338
rect 10769 3738 10897 4338
rect 10925 3738 10981 4338
rect 11081 3738 11131 4338
rect 12916 4209 12966 4264
rect 531 2658 584 2808
rect 534 2208 584 2658
rect 704 2208 760 2808
rect 880 2208 936 2808
rect 1056 2208 1112 2808
rect 1232 2208 1282 2808
rect 1348 2208 1398 2808
rect 1518 2208 1574 2808
rect 1694 2208 1750 2808
rect 1870 2208 1920 2808
rect 2191 2608 2371 2808
rect 2427 2608 2607 2808
rect 4161 2608 4341 2808
rect 4397 2608 4577 2808
rect 2427 2473 2607 2510
rect 4161 2473 4341 2510
rect 4848 2208 4898 2808
rect 5018 2208 5074 2808
rect 5194 2208 5250 2808
rect 5370 2208 5420 2808
rect 5502 2208 5552 2808
rect 5672 2208 5728 2808
rect 5848 2208 5904 2808
rect 6024 2208 6074 2808
rect 6345 2608 6525 2808
rect 6581 2608 6761 2808
rect 8315 2608 8495 2808
rect 8551 2608 8731 2808
rect 6581 2473 6761 2510
rect 8315 2473 8495 2510
rect 9002 2208 9052 2808
rect 9172 2208 9228 2808
rect 9348 2208 9404 2808
rect 9524 2208 9574 2808
rect 9656 2208 9706 2808
rect 9826 2208 9882 2808
rect 10002 2208 10058 2808
rect 10178 2208 10228 2808
rect 10499 2608 10679 2808
rect 10735 2608 10915 2808
rect 12469 2608 12649 2808
rect 12705 2608 12885 2808
rect 10735 2473 10915 2510
rect 12469 2473 12649 2510
rect 13156 2208 13206 2808
rect 13326 2208 13382 2808
rect 13502 2208 13558 2808
rect 13678 2208 13728 2808
rect 13909 1810 13933 1834
rect 14330 1810 14354 1834
rect 13933 1786 13957 1801
rect 14306 1786 14330 1801
rect 13737 1630 13761 1654
rect 13762 1606 13785 1630
rect 157 792 207 1392
rect 327 792 383 1392
rect 503 792 553 1392
rect 2046 1000 2096 1600
rect 2216 1000 2266 1600
rect 2642 995 2692 1595
rect 2812 995 2868 1595
rect 2988 1348 3038 1595
rect 3101 1445 3113 1595
rect 3727 1445 3780 1595
rect 3730 1348 3780 1445
rect 2988 1276 3041 1348
rect 2988 995 3038 1276
rect 3101 1126 3113 1276
rect 3727 1126 3780 1348
rect 3730 995 3780 1126
rect 3900 995 3956 1595
rect 4076 995 4126 1595
rect 4502 1000 4552 1600
rect 4672 1000 4722 1600
rect 6200 1000 6250 1600
rect 6370 1000 6420 1600
rect 6796 995 6846 1595
rect 6966 995 7022 1595
rect 7142 1348 7192 1595
rect 7255 1445 7267 1595
rect 7881 1445 7934 1595
rect 7884 1348 7934 1445
rect 7142 1276 7195 1348
rect 7142 995 7192 1276
rect 7255 1126 7267 1276
rect 7881 1126 7934 1348
rect 7884 995 7934 1126
rect 8054 995 8110 1595
rect 8230 995 8280 1595
rect 8656 1000 8706 1600
rect 8826 1000 8876 1600
rect 10354 1000 10404 1600
rect 10524 1000 10574 1600
rect 10950 995 11000 1595
rect 11120 995 11176 1595
rect 11296 1348 11346 1595
rect 11409 1445 11421 1595
rect 12035 1445 12088 1595
rect 12038 1348 12088 1445
rect 11296 1276 11349 1348
rect 11296 995 11346 1276
rect 11409 1126 11421 1276
rect 12035 1126 12088 1348
rect 12038 995 12088 1126
rect 12208 995 12264 1595
rect 12384 995 12434 1595
rect 12810 1000 12860 1600
rect 12980 1000 13030 1600
rect 13957 1542 13991 1566
rect 14027 1542 14061 1566
rect 14097 1542 14131 1566
rect 14167 1542 14201 1566
rect 14237 1542 14271 1566
rect 14307 1542 14330 1566
rect 13762 1508 13785 1532
rect 13737 1484 13761 1508
rect 1585 673 1619 697
rect 1653 673 1687 697
rect 1721 673 1755 697
rect 1789 673 1823 697
rect 1857 673 1891 697
rect 1925 673 1959 697
rect 1993 673 2027 697
rect 2061 673 2095 697
rect 2129 673 2163 697
rect 2197 673 2231 697
rect 2265 673 2299 697
rect 2333 673 2367 697
rect 2401 673 2435 697
rect 2469 673 2503 697
rect 2537 673 2571 697
rect 2605 673 2639 697
rect 2673 673 2707 697
rect 2741 673 2775 697
rect 2809 673 2843 697
rect 2877 673 2911 697
rect 2945 673 2979 697
rect 3013 673 3047 697
rect 3081 673 3115 697
rect 3149 673 3183 697
rect 3217 673 3251 697
rect 3285 673 3319 697
rect 3353 673 3387 697
rect 3421 673 3455 697
rect 3489 673 3523 697
rect 3557 673 3591 697
rect 3625 673 3659 697
rect 3693 673 3727 697
rect 3761 673 3795 697
rect 3829 673 3863 697
rect 3897 673 3931 697
rect 3965 673 3999 697
rect 4033 673 4067 697
rect 4101 673 4135 697
rect 4169 673 4203 697
rect 4237 673 4271 697
rect 4305 673 4339 697
rect 4373 673 4407 697
rect 4441 673 4475 697
rect 4509 673 4543 697
rect 4577 673 4611 697
rect 4645 673 4679 697
rect 4713 673 4747 697
rect 4781 673 4815 697
rect 4849 673 4883 697
rect 4917 673 4951 697
rect 4985 673 5019 697
rect 5053 673 5087 697
rect 5121 673 5155 697
rect 5189 673 5223 697
rect 5257 673 5291 697
rect 5325 673 5359 697
rect 5393 673 5427 697
rect 5461 673 5495 697
rect 5529 673 5563 697
rect 5597 673 5631 697
rect 5665 673 5699 697
rect 5733 673 5767 697
rect 5801 673 5835 697
rect 5869 673 5903 697
rect 5937 673 5971 697
rect 6005 673 6039 697
rect 6073 673 6107 697
rect 6141 673 6175 697
rect 6209 673 6243 697
rect 6277 673 6311 697
rect 6345 673 6379 697
rect 6413 673 6447 697
rect 6481 673 6515 697
rect 6549 673 6583 697
rect 6617 673 6651 697
rect 6685 673 6719 697
rect 6753 673 6787 697
rect 6821 673 6855 697
rect 6889 673 6923 697
rect 6957 673 6991 697
rect 7025 673 7059 697
rect 7093 673 7127 697
rect 7161 673 7195 697
rect 7229 673 7263 697
rect 7297 673 7331 697
rect 7365 673 7399 697
rect 7433 673 7467 697
rect 7501 673 7535 697
rect 7569 673 7603 697
rect 7637 673 7671 697
rect 7705 673 7739 697
rect 7773 673 7807 697
rect 7841 673 7875 697
rect 7909 673 7943 697
rect 7977 673 8011 697
rect 8045 673 8079 697
rect 8113 673 8147 697
rect 8181 673 8215 697
rect 8249 673 8283 697
rect 8317 673 8351 697
rect 8385 673 8419 697
rect 8453 673 8487 697
rect 8521 673 8555 697
rect 8589 673 8623 697
rect 8657 673 8691 697
rect 8725 673 8759 697
rect 8793 673 8827 697
rect 8861 673 8895 697
rect 8929 673 8963 697
rect 9063 673 9097 697
rect 9131 673 9165 697
rect 9199 673 9233 697
rect 9267 673 9301 697
rect 9335 673 9369 697
rect 9403 673 9437 697
rect 9471 673 9505 697
rect 9539 673 9573 697
rect 9607 673 9641 697
rect 9675 673 9709 697
rect 9743 673 9777 697
rect 9811 673 9845 697
rect 9879 673 9913 697
rect 9947 673 9981 697
rect 10015 673 10049 697
rect 10083 673 10117 697
rect 10151 673 10185 697
rect 10219 673 10253 697
rect 10287 673 10321 697
rect 10355 673 10389 697
rect 10423 673 10457 697
rect 10491 673 10525 697
rect 10559 673 10593 697
rect 10627 673 10661 697
rect 10695 673 10729 697
rect 10763 673 10797 697
rect 10831 673 10865 697
rect 10899 673 10933 697
rect 10967 673 11001 697
rect 11035 673 11069 697
rect 11103 673 11137 697
rect 11171 673 11205 697
rect 11239 673 11273 697
rect 11307 673 11341 697
rect 11375 673 11409 697
rect 11443 673 11477 697
rect 11511 673 11545 697
rect 11579 673 11613 697
rect 11647 673 11681 697
rect 11715 673 11749 697
rect 11783 673 11817 697
rect 11851 673 11885 697
rect 11919 673 11953 697
rect 11987 673 12021 697
rect 12055 673 12089 697
rect 12123 673 12157 697
rect 9013 647 9039 673
<< metal1 >>
rect 12486 -407 12538 -351
<< metal2 >>
rect 7956 15977 8019 15991
rect 7956 15927 7969 15977
tri 7969 15927 8019 15977 nw
rect 675 -407 721 -361
rect 1084 -407 1130 -328
rect 1226 -407 1278 -355
rect 2551 -407 2603 -363
rect 3262 -407 3314 -306
rect 4471 -407 4523 -340
rect 5320 -407 5372 -379
rect 5698 -407 5750 -355
rect 6150 -407 6202 -351
rect 6363 -407 6415 -363
rect 7092 -407 7144 -351
rect 7678 -407 7730 -318
rect 9049 -407 9101 -355
rect 9971 -407 10023 -355
rect 13367 -407 13419 -355
rect 13655 -407 13785 -363
rect 15256 -407 15384 -363
rect 15522 -407 15574 -363
rect 15741 -407 15781 -363
rect 15943 -407 15983 -215
<< metal3 >>
rect 80 -407 204 -244
rect 9173 -407 9239 -355
rect 12564 -407 12778 -260
rect 15716 -407 15782 -254
rect 15848 -407 15914 -244
<< metal4 >>
rect 0 34750 254 39593
rect 15746 34750 16000 39593
rect 0 13600 254 18593
rect 15746 13600 16000 18593
rect 0 12410 254 13300
rect 15746 12410 16000 13300
rect 0 11240 254 12130
rect 15746 11240 16000 12130
rect 0 10874 254 10940
rect 15746 10874 16000 10940
rect 0 10218 100 10814
rect 15746 10218 15846 10814
rect 0 9922 254 10158
rect 15746 9922 16000 10158
rect 0 9266 116 9862
rect 15746 9266 15862 9862
rect 0 9140 254 9206
rect 15746 9140 16000 9206
rect 0 7910 254 8840
rect 15746 7910 16000 8840
rect 0 6940 254 7630
rect 15746 6940 16000 7630
rect 0 5970 254 6660
rect 15746 5970 16000 6660
rect 0 4760 254 5690
rect 15746 4760 16000 5690
rect 0 3550 254 4480
rect 15746 3550 16000 4480
rect 0 2580 254 3270
rect 15746 2580 16000 3270
rect 0 1370 254 2300
rect 15746 1370 16000 2300
rect 0 0 254 1090
rect 15746 0 16000 1090
<< metal5 >>
rect 0 34750 254 39593
rect 15746 34750 16000 39593
rect 6423 24687 10731 28996
rect 0 13600 254 18590
rect 15746 13600 16000 18590
rect 0 12430 254 13280
rect 15746 12430 16000 13280
rect 0 11260 254 12110
rect 15746 11260 16000 12110
rect 0 9140 254 10940
rect 15746 9140 16000 10940
rect 0 7930 254 8820
rect 15746 7930 16000 8820
rect 0 6960 254 7610
rect 15746 6960 16000 7610
rect 0 5990 254 6640
rect 15746 5990 16000 6640
rect 0 4780 254 5670
rect 15746 4780 16000 5670
rect 0 3570 254 4460
rect 15746 3570 16000 4460
rect 0 2600 254 3250
rect 15746 2600 16000 3250
rect 0 1390 254 2280
rect 15746 1390 16000 2280
rect 0 20 254 1070
rect 15746 20 16000 1070
use sky130_fd_io__top_gpiov2  sky130_fd_io__top_gpiov2_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602555073
transform 1 0 0 0 1 -407
box -143 -136 16134 40000
use sky130_fd_io__overlay_gpiov2  sky130_fd_io__overlay_gpiov2_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602555073
transform 1 0 0 0 1 -407
box 0 407 16000 40000
<< labels >>
flabel metal4 s 127 37925 127 37925 3 FreeSans 520 0 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal5 s 0 13600 254 18590 3 FreeSans 520 0 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal5 s 0 7930 254 8820 3 FreeSans 520 0 0 0 VSSD
port 34 nsew ground bidirectional
flabel metal5 s 0 11260 254 12110 3 FreeSans 520 0 0 0 VSSIO_Q
port 36 nsew ground bidirectional
flabel metal5 s 0 5990 254 6640 3 FreeSans 520 0 0 0 VSWITCH
port 37 nsew power bidirectional
flabel metal5 s 0 4780 254 5670 3 FreeSans 520 0 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal5 s 0 2600 193 3250 3 FreeSans 520 0 0 0 VDDA
port 30 nsew power bidirectional
flabel metal5 s 0 3570 254 4460 3 FreeSans 520 0 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal5 s 0 1390 254 2280 3 FreeSans 520 0 0 0 VCCD
port 28 nsew power bidirectional
flabel metal5 s 0 12430 254 13280 3 FreeSans 520 0 0 0 VDDIO_Q
port 32 nsew power bidirectional
flabel metal5 s 0 9140 254 10940 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal5 s 0 6961 254 7610 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal5 s 0 20 254 1070 3 FreeSans 520 0 0 0 VCCHIB
port 29 nsew power bidirectional
flabel metal4 s 0 34750 254 39593 3 FreeSans 520 0 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal4 s 0 3550 254 4480 3 FreeSans 520 0 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal4 s 0 12410 254 13300 3 FreeSans 520 0 0 0 VDDIO_Q
port 32 nsew power bidirectional
flabel metal4 s 0 13600 254 18593 3 FreeSans 520 0 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal4 s 0 1370 254 2300 3 FreeSans 520 0 0 0 VCCD
port 28 nsew power bidirectional
flabel metal4 s 0 9140 254 9206 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 0 5970 254 6660 3 FreeSans 520 0 0 0 VSWITCH
port 37 nsew power bidirectional
flabel metal4 s 0 9922 254 10158 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 0 11240 254 12130 3 FreeSans 520 0 0 0 VSSIO_Q
port 36 nsew ground bidirectional
flabel metal4 s 0 4760 254 5690 3 FreeSans 520 0 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal4 s 0 2580 193 3270 3 FreeSans 520 0 0 0 VDDA
port 30 nsew power bidirectional
flabel metal4 s 0 10218 254 10814 3 FreeSans 520 0 0 0 AMUXBUS_A
port 0 nsew signal bidirectional
flabel metal4 s 0 10874 254 10940 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 0 6940 254 7630 3 FreeSans 520 0 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 0 7910 254 8840 3 FreeSans 520 0 0 0 VSSD
port 34 nsew ground bidirectional
flabel metal4 s 0 9266 254 9862 3 FreeSans 520 0 0 0 AMUXBUS_B
port 1 nsew signal bidirectional
flabel metal4 s 0 0 254 1090 3 FreeSans 520 0 0 0 VCCHIB
port 29 nsew power bidirectional
flabel metal4 s 15873 37925 15873 37925 3 FreeSans 520 180 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal5 s 15746 9140 16000 10940 3 FreeSans 520 180 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal5 s 15807 2600 16000 3250 3 FreeSans 520 180 0 0 VDDA
port 30 nsew power bidirectional
flabel metal5 s 15746 7930 16000 8820 3 FreeSans 520 180 0 0 VSSD
port 34 nsew ground bidirectional
flabel metal5 s 15746 11260 16000 12110 3 FreeSans 520 180 0 0 VSSIO_Q
port 36 nsew ground bidirectional
flabel metal5 s 15746 4780 16000 5670 3 FreeSans 520 180 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal5 s 15746 5990 16000 6640 3 FreeSans 520 180 0 0 VSWITCH
port 37 nsew power bidirectional
flabel metal5 s 15746 6961 16000 7610 3 FreeSans 520 180 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal5 s 15746 1390 16000 2280 3 FreeSans 520 180 0 0 VCCD
port 28 nsew power bidirectional
flabel metal5 s 15746 12430 16000 13280 3 FreeSans 520 180 0 0 VDDIO_Q
port 32 nsew power bidirectional
flabel metal5 s 15746 13600 16000 18590 3 FreeSans 520 180 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal5 s 15746 20 16000 1070 3 FreeSans 520 180 0 0 VCCHIB
port 29 nsew power bidirectional
flabel metal5 s 15746 3570 16000 4460 3 FreeSans 520 180 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal4 s 15746 7910 16000 8840 3 FreeSans 520 180 0 0 VSSD
port 34 nsew ground bidirectional
flabel metal4 s 15807 2580 16000 3270 3 FreeSans 520 180 0 0 VDDA
port 30 nsew power bidirectional
flabel metal4 s 15746 11240 16000 12130 3 FreeSans 520 180 0 0 VSSIO_Q
port 36 nsew ground bidirectional
flabel metal4 s 15746 4760 16000 5690 3 FreeSans 520 180 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal4 s 15746 5970 16000 6660 3 FreeSans 520 180 0 0 VSWITCH
port 37 nsew power bidirectional
flabel metal4 s 15746 9922 16000 10158 3 FreeSans 520 180 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 15746 10874 16000 10940 3 FreeSans 520 180 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 15746 3550 16000 4480 3 FreeSans 520 180 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal4 s 15746 9140 16000 9206 3 FreeSans 520 180 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 15746 6940 16000 7630 3 FreeSans 520 180 0 0 VSSA
port 33 nsew ground bidirectional
flabel metal4 s 15746 12410 16000 13300 3 FreeSans 520 180 0 0 VDDIO_Q
port 32 nsew power bidirectional
flabel metal4 s 15746 1370 16000 2300 3 FreeSans 520 180 0 0 VCCD
port 28 nsew power bidirectional
flabel metal4 s 15746 9266 16000 9862 3 FreeSans 520 180 0 0 AMUXBUS_B
port 1 nsew signal bidirectional
flabel metal4 s 15746 34750 16000 39593 3 FreeSans 520 180 0 0 VSSIO
port 35 nsew ground bidirectional
flabel metal4 s 15746 10218 16000 10814 3 FreeSans 520 180 0 0 AMUXBUS_A
port 0 nse signal bidirectional
flabel metal4 s 15746 13600 16000 18593 3 FreeSans 520 180 0 0 VDDIO
port 31 nsew power bidirectional
flabel metal4 s 15746 0 16000 1090 3 FreeSans 520 180 0 0 VCCHIB
port 29 nsew power bidirectional
flabel metal5 s 6423 24687 10731 28996 0 FreeSans 1600 0 0 0 PAD
port 21 nsew signal bidirectional
flabel metal3 s 80 -407 204 -244 0 FreeSans 640 0 0 0 IN_H
port 17 nsew signal output
flabel metal2 s 675 -407 721 -361 0 FreeSans 400 270 0 0 OE_N
port 19 nsew signal input
flabel metal2 s 1084 -407 1130 -328 0 FreeSans 400 270 0 0 IB_MODE_SEL
port 15 nsew signal input
flabel metal2 s 1226 -407 1278 -355 0 FreeSans 400 270 0 0 VTRIP_SEL
port 38 nsew signal input
flabel metal2 s 2551 -407 2603 -363 0 FreeSans 400 270 0 0 ENABLE_VDDA_H
port 10 nsew signal input
flabel metal2 s 3262 -407 3314 -306 0 FreeSans 400 270 0 0 ENABLE_VSWITCH_H
port 12 nsew signal input
flabel metal2 s 4471 -407 4523 -340 0 FreeSans 400 0 0 0 OUT
port 20 nsew signal input
flabel metal2 s 5320 -407 5372 -379 0 FreeSans 400 270 0 0 HLD_OVR
port 14 nsew signal input
flabel metal2 s 5698 -407 5750 -355 0 FreeSans 400 270 0 0 DM[2]
port 5 nsew signal input
flabel metal2 s 6150 -407 6202 -351 0 FreeSans 400 270 0 0 ANALOG_SEL
port 4 nsew signal input
flabel metal2 s 6363 -407 6415 -363 0 FreeSans 400 270 0 0 HLD_H_N
port 13 nsew signal input
flabel metal2 s 7092 -407 7144 -351 0 FreeSans 400 270 0 0 ENABLE_H
port 8 nsew signal input
flabel metal2 s 7678 -407 7730 -318 0 FreeSans 400 270 0 0 ENABLE_INP_H
port 9 nsew signal input
flabel metal2 s 9049 -407 9101 -355 0 FreeSans 400 270 0 0 INP_DIS
port 18 nsew signal input
flabel metal3 s 9173 -407 9239 -355 0 FreeSans 400 270 0 0 ANALOG_POL
port 3 nsew signal input
flabel metal2 s 9971 -407 10023 -355 0 FreeSans 400 270 0 0 DM[0]
port 7 nsew signal input
flabel metal1 s 12486 -407 12538 -351 0 FreeSans 400 270 0 0 ANALOG_EN
port 2 nsew signal input
flabel metal2 s 13367 -407 13419 -355 0 FreeSans 400 270 0 0 DM[1]
port 6 nsew signal input
flabel metal2 s 15522 -407 15574 -363 0 FreeSans 400 270 0 0 SLOW
port 25 nsew signal input
flabel metal3 s 15848 -407 15914 -244 0 FreeSans 400 270 0 0 IN
port 16 nsew signal output
flabel metal3 s 12564 -407 12778 -260 0 FreeSans 400 270 0 0 PAD_A_NOESD_H
port 24 nsew signal bidirectional
flabel metal2 s 13655 -407 13785 -363 0 FreeSans 400 270 0 0 PAD_A_ESD_1_H
port 23 nsew signal bidirectional
flabel metal2 s 15256 -407 15384 -363 0 FreeSans 400 270 0 0 PAD_A_ESD_0_H
port 22 nsew signal bidirectional
flabel metal2 s 15943 -407 15983 -215 0 FreeSans 400 270 0 0 TIE_LO_ESD
port 27 nsew signal output
flabel metal2 s 15741 -407 15781 -363 0 FreeSans 400 270 0 0 TIE_HI_ESD
port 26 nsew signal output
flabel metal3 s 15716 -407 15782 -254 0 FreeSans 400 270 0 0 ENABLE_VDDIO
port 11 nsew signal input
<< properties >>
string LEFclass PAD INOUT
string FIXED_BBOX 0 0 16000 39593
<< end >>
