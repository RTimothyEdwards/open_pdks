magic
tech sky130A
magscale 1 2
timestamp 1602972891
<< error_p >>
rect 1419 2270 1664 2276
rect 2097 2235 2343 2239
rect 2096 2207 2342 2211
rect 3193 2209 3227 2243
rect 3634 2215 3671 2255
rect 2673 2183 2679 2189
rect 2731 2183 2737 2189
rect 2679 2177 2685 2180
rect 2725 2177 2731 2180
rect 1407 1398 1449 1423
rect 1407 1342 1449 1367
rect 3303 1040 3320 1367
<< metal1 >>
rect 2679 2235 2731 2308
rect 2679 2180 2731 2183
<< via1 >>
rect 2679 2183 2731 2235
<< metal2 >>
rect 1419 2248 1664 2270
rect 2097 2235 2343 2272
rect 3589 2255 3716 2300
rect 2096 2174 2342 2211
rect 2670 2183 2679 2235
rect 2731 2183 2787 2235
rect 3193 2209 3227 2243
rect 3589 2215 3634 2255
rect 3671 2215 3716 2255
rect 3589 2170 3716 2215
rect 1449 1433 2149 1583
rect 1407 1398 2149 1433
rect 1449 1367 2149 1398
rect 1407 1332 2149 1367
rect 1449 883 2149 1332
rect 2564 866 3264 1566
rect 3303 1040 3332 1367
<< labels >>
flabel comment s 500 1677 500 1677 0 FreeSans 560 0 0 0 Not implemented
flabel comment s 493 2348 493 2348 0 FreeSans 800 0 0 0 Met2 (m2)
flabel comment s 568 1459 568 1459 0 FreeSans 560 0 0 0 m2.4a
flabel comment s 1549 2081 1549 2081 0 FreeSans 560 0 0 0 m2.1
flabel comment s 2260 2050 2260 2050 0 FreeSans 560 0 0 0 m2.2
flabel comment s 1821 811 1821 811 0 FreeSans 560 0 0 0 m2.3a
flabel comment s 2974 811 2974 811 0 FreeSans 560 0 0 0 m2.3b
flabel comment s 505 2126 505 2126 0 FreeSans 560 0 0 0 Correct by design
flabel comment s 530 2005 530 2005 0 FreeSans 560 0 0 0 m2.4
flabel comment s 2740 2110 2740 2110 0 FreeSans 560 0 0 0 m2.5
flabel comment s 3238 2101 3238 2101 0 FreeSans 560 0 0 0 m2.6
flabel comment s 3630 2099 3630 2099 0 FreeSans 560 0 0 0 m2.7
<< end >>
