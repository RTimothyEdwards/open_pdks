VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_io__com_bus_slice_10um
  CLASS PAD SPACER ;
  FOREIGN sky130_ef_io__com_bus_slice_10um ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 10.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 10.000 49.310 ;
    END
  END AMUXBUS_B
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 10.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 10.000 46.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.800 10.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 10.000 38.150 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 10.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 10.000 16.350 ;
    END
  END VDDA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 10.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 10.000 33.300 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 10.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 10.000 66.500 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 10.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 10.000 5.450 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 10.000 92.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 10.000 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 10.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 10.000 22.400 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 10.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 10.000 11.500 ;
    END
  END VCCD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 10.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 10.000 28.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.750 10.000 197.965 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 10.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 10.000 44.200 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 10.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 10.000 60.650 ;
    END
  END VSSIO_Q
  OBS
      LAYER met4 ;
        RECT 0.000 173.75 10.000 197.965 ;
        RECT 0.000 66.900 10.000 67.600 ;
        RECT 0.000 61.050 10.000 61.650 ;
        RECT 0.000 55.100 10.000 55.800 ;
        RECT 0.000 49.610 10.000 50.790 ;
  END
END sky130_ef_io__com_bus_slice_10um
END LIBRARY

