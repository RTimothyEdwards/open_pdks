VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_io__gpiov2_pad
  CLASS PAD INOUT ;
  FOREIGN sky130_ef_io__gpiov2_pad ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 197.965 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.090 36.440 54.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.760 51.090 80.000 54.070 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.330 52.145 49.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.465 46.330 80.000 49.310 ;
    END
  END AMUXBUS_B
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430 -2.035 62.690 -0.730 ;
    END
  END ANALOG_EN
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865 -2.035 46.195 34.770 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.750 -2.035 31.010 0.230 ;
    END
  END ANALOG_SEL
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490 -2.035 28.750 2.035 ;
    END
  END DM[2]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.835 -2.035 67.095 -0.840 ;
    END
  END DM[1]
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.855 -2.035 50.115 -1.490 ;
    END
  END DM[0]
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.460 -2.035 35.720 -0.485 ;
    END
  END ENABLE_H
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390 -2.035 38.650 1.055 ;
    END
  END ENABLE_INP_H
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.755 -2.035 13.015 3.315 ;
    END
  END ENABLE_VDDA_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580 -2.035 78.910 182.740 ;
    END
  END ENABLE_VDDIO
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.310 -2.035 16.570 0.285 ;
    END
  END ENABLE_VSWITCH_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815 -2.035 32.075 1.305 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600 -2.035 26.860 0.670 ;
    END
  END HLD_OVR
  PIN IB_MODE_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420 -2.035 5.650 2.440 ;
    END
  END IB_MODE_SEL
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240 -2.035 79.570 187.525 ;
    END
  END IN
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400 -2.035 1.020 176.450 ;
    END
  END IN_H
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245 -2.035 45.505 3.055 ;
    END
  END INP_DIS
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375 -2.035 3.605 2.440 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355 -2.035 22.615 4.390 ;
    END
  END OUT
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.200 102.525 73.800 164.975 ;
    END
  END PAD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280 -2.035 76.920 0.020 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275 -2.035 68.925 0.235 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.820 -2.035 63.890 7.670 ;
    END
  END PAD_A_NOESD_H
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.610 -2.035 77.870 -0.850 ;
    END
  END SLOW
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.705 -2.035 78.905 -0.820 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715 -2.035 79.915 175.835 ;
    END
  END TIE_LO_ESD
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.950 1.270 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.850 1.270 11.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 6.950 80.000 11.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 6.850 80.000 11.500 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.100 1.270 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.000 1.270 5.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 0.100 80.000 5.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 0.000 80.000 5.450 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.000 0.965 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.900 0.965 16.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.970 13.000 80.000 16.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 12.900 80.000 16.350 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.000 1.270 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.850 1.270 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.750 1.270 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.000 1.270 92.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 68.000 80.000 92.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 17.850 80.000 22.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 17.750 80.000 22.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 68.000 80.000 92.965 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.150 1.270 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.050 1.270 66.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 62.150 80.000 66.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 62.050 80.000 66.500 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.700 1.270 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.805 1.270 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.700 2.610 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.610 1.270 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.370 2.610 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.700 1.270 38.150 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 45.700 80.000 54.700 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 34.805 80.000 38.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 49.610 80.000 50.790 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 54.370 80.000 54.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 45.700 80.000 46.030 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 34.700 80.000 38.150 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.650 1.270 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.550 1.270 44.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 39.650 80.000 44.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 39.550 80.000 44.200 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 0.810 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.900 1.270 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.750 1.270 197.965 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.800 1.270 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 173.750 80.000 197.965 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 23.900 80.000 28.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 23.800 80.000 28.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 173.750 80.000 197.965 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.300 1.270 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.200 1.270 60.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 56.300 80.000 60.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 56.200 80.000 60.650 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.950 1.270 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.850 1.270 33.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 29.950 80.000 33.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 29.850 80.000 33.300 ;
    END
  END VSWITCH
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130 -2.035 6.390 -0.485 ;
    END
  END VTRIP_SEL
  OBS
      LAYER nwell ;
        RECT -0.415 171.510 80.435 176.940 ;
        RECT -0.415 168.440 7.515 171.510 ;
        RECT 66.970 168.440 80.435 171.510 ;
        RECT -0.415 168.195 80.435 168.440 ;
        RECT -0.415 166.480 80.440 168.195 ;
        RECT -0.415 144.655 6.385 166.480 ;
        RECT 78.630 144.655 80.440 166.480 ;
        RECT -0.415 142.845 80.440 144.655 ;
      LAYER pwell ;
        RECT -0.160 138.780 80.160 142.400 ;
      LAYER nwell ;
        RECT 46.040 138.345 80.440 138.350 ;
        RECT -0.415 128.630 80.440 138.345 ;
      LAYER pwell ;
        RECT -0.085 127.150 40.115 128.190 ;
        RECT 67.040 127.150 80.160 128.190 ;
        RECT -0.085 123.230 80.160 127.150 ;
        RECT -0.085 101.385 5.605 123.230 ;
        RECT 77.995 101.385 80.160 123.230 ;
        RECT -0.085 100.060 80.160 101.385 ;
        RECT -0.085 94.090 5.085 100.060 ;
        RECT 39.515 98.915 80.160 100.060 ;
        RECT 53.010 97.615 80.160 98.915 ;
        RECT 76.900 95.820 80.160 97.615 ;
        RECT 39.515 94.090 80.160 95.820 ;
        RECT -0.085 94.070 80.160 94.090 ;
        RECT -0.085 93.095 45.710 94.070 ;
        RECT -0.085 93.050 46.460 93.095 ;
        RECT -0.085 91.030 9.170 93.050 ;
      LAYER nwell ;
        RECT 46.940 92.210 80.670 93.130 ;
        RECT 62.650 91.700 80.670 92.210 ;
        RECT -0.415 89.785 2.795 90.365 ;
        RECT -0.415 86.450 5.975 89.785 ;
        RECT -0.120 86.245 5.975 86.450 ;
        RECT -0.120 85.705 8.420 86.245 ;
        RECT -0.120 84.625 8.495 85.705 ;
        RECT -0.120 83.545 4.530 84.625 ;
        RECT 79.240 82.310 80.670 91.700 ;
        RECT 46.940 81.130 80.670 82.310 ;
        RECT -0.715 77.770 24.815 79.200 ;
        RECT -0.715 60.305 0.715 77.770 ;
        RECT 79.240 71.740 80.670 81.130 ;
        RECT 62.650 71.230 80.670 71.740 ;
        RECT 46.940 70.560 80.670 71.230 ;
        RECT 79.125 64.010 80.670 70.560 ;
        RECT 70.335 63.160 80.670 64.010 ;
        RECT -0.715 58.985 3.810 60.305 ;
        RECT -0.715 58.735 13.535 58.985 ;
        RECT -0.715 58.145 10.460 58.735 ;
        RECT -0.715 55.985 0.715 58.145 ;
        RECT -0.715 54.555 23.515 55.985 ;
        RECT 79.125 50.015 80.670 63.160 ;
        RECT 70.335 48.585 80.670 50.015 ;
        RECT 48.915 32.230 80.450 34.020 ;
        RECT 58.275 30.375 80.450 32.230 ;
        RECT 64.830 27.750 80.450 30.375 ;
        RECT 64.830 21.045 80.450 23.310 ;
        RECT 4.580 17.120 80.450 21.045 ;
        RECT -0.415 3.630 3.110 7.290 ;
        RECT 0.000 -2.035 61.490 1.465 ;
        RECT 64.030 -0.145 65.390 2.135 ;
      LAYER pwell ;
        RECT 64.375 -1.785 66.075 -1.035 ;
      LAYER li1 ;
        RECT 0.000 176.610 80.000 197.670 ;
        RECT -0.085 168.055 80.105 176.610 ;
        RECT -0.115 143.180 80.105 168.055 ;
        RECT -0.115 143.120 80.000 143.180 ;
        RECT 0.000 142.400 80.000 143.120 ;
        RECT -0.160 138.780 80.160 142.400 ;
        RECT 0.000 138.115 80.000 138.780 ;
        RECT -0.115 138.020 80.000 138.115 ;
        RECT -0.115 129.240 80.085 138.020 ;
        RECT -0.085 128.960 80.085 129.240 ;
        RECT 0.000 128.190 80.000 128.960 ;
        RECT -0.085 128.185 80.160 128.190 ;
        RECT -0.115 94.070 80.160 128.185 ;
        RECT -0.115 93.860 80.000 94.070 ;
        RECT -0.085 92.545 80.000 93.860 ;
        RECT -0.085 91.030 80.085 92.545 ;
        RECT 0.000 90.035 80.085 91.030 ;
        RECT -0.085 86.780 80.085 90.035 ;
        RECT 0.000 78.570 80.085 86.780 ;
        RECT -0.085 55.185 80.085 78.570 ;
        RECT 0.000 49.215 80.085 55.185 ;
        RECT 0.000 33.690 80.000 49.215 ;
        RECT 0.000 28.080 80.120 33.690 ;
        RECT 0.000 22.980 80.000 28.080 ;
        RECT 0.000 17.450 80.120 22.980 ;
        RECT 0.000 6.960 80.000 17.450 ;
        RECT -0.085 3.960 80.000 6.960 ;
        RECT 0.000 0.000 80.000 3.960 ;
        RECT 0.705 -0.100 0.875 0.000 ;
        RECT 0.705 -0.520 1.625 -0.100 ;
        RECT 2.090 -0.485 2.420 0.000 ;
        RECT 0.705 -1.500 0.875 -0.830 ;
        RECT 1.485 -0.860 1.655 -0.830 ;
        RECT 1.485 -1.390 1.660 -0.860 ;
        RECT 2.590 -1.345 2.760 0.000 ;
        RECT 3.470 -1.195 3.640 0.000 ;
        RECT 3.830 -0.080 4.160 0.000 ;
        RECT 4.350 -1.345 4.520 0.000 ;
        RECT 5.230 -1.195 5.400 0.000 ;
        RECT 6.110 -1.345 6.280 0.000 ;
        RECT 6.730 -1.345 6.900 0.000 ;
        RECT 7.610 -1.205 7.780 0.000 ;
        RECT 8.490 -1.345 8.660 0.000 ;
        RECT 9.370 -1.205 9.540 0.000 ;
        RECT 10.250 -1.345 10.420 0.000 ;
        RECT 10.615 -0.055 10.945 0.000 ;
        RECT 11.130 -1.205 11.300 0.000 ;
        RECT 11.750 -1.345 11.920 0.000 ;
        RECT 12.630 -1.205 12.800 0.000 ;
        RECT 13.510 -1.345 13.680 0.000 ;
        RECT 14.390 -1.205 14.560 0.000 ;
        RECT 15.270 -1.345 15.440 0.000 ;
        RECT 16.150 -1.205 16.320 0.000 ;
        RECT 17.030 -1.345 17.200 0.000 ;
        RECT 17.910 -1.205 18.080 0.000 ;
        RECT 18.790 -1.345 18.960 0.000 ;
        RECT 19.670 -1.205 19.840 0.000 ;
        RECT 20.550 -1.345 20.720 0.000 ;
        RECT 21.430 -1.205 21.600 0.000 ;
        RECT 22.310 -1.345 22.480 0.000 ;
        RECT 23.190 -1.205 23.360 0.000 ;
        RECT 24.070 -1.345 24.240 0.000 ;
        RECT 24.950 -1.205 25.120 0.000 ;
        RECT 25.830 -1.345 26.000 0.000 ;
        RECT 26.710 -1.205 26.880 0.000 ;
        RECT 27.590 -1.345 27.760 0.000 ;
        RECT 28.470 -1.205 28.640 0.000 ;
        RECT 29.350 -1.345 29.520 0.000 ;
        RECT 29.965 -0.050 30.495 0.000 ;
        RECT 29.970 -1.205 30.140 -0.050 ;
        RECT 30.850 -1.345 31.020 0.000 ;
        RECT 31.470 -1.345 31.640 0.000 ;
        RECT 32.350 -1.205 32.520 0.000 ;
        RECT 33.230 -1.345 33.400 0.000 ;
        RECT 34.110 -0.265 34.285 0.000 ;
        RECT 34.110 -1.205 34.280 -0.265 ;
        RECT 37.990 -1.345 38.160 0.000 ;
        RECT 38.870 -1.205 39.040 0.000 ;
        RECT 39.750 -1.345 39.920 0.000 ;
        RECT 40.630 -1.205 40.800 0.000 ;
        RECT 41.250 -1.345 41.420 0.000 ;
        RECT 42.130 -1.195 42.300 0.000 ;
        RECT 43.010 -1.345 43.180 0.000 ;
        RECT 45.290 -0.410 45.460 0.000 ;
        RECT 45.110 -0.580 45.640 -0.410 ;
        RECT 45.290 -1.205 45.460 -0.580 ;
        RECT 46.170 -1.345 46.340 0.000 ;
        RECT 47.050 -1.195 47.220 0.000 ;
        RECT 47.930 -1.345 48.100 0.000 ;
        RECT 48.495 -1.345 48.665 0.000 ;
        RECT 49.375 -1.205 49.545 0.000 ;
        RECT 50.255 -1.345 50.425 0.000 ;
        RECT 51.135 -1.205 51.305 0.000 ;
        RECT 52.015 -1.345 52.185 0.000 ;
        RECT 52.640 -1.205 52.810 0.000 ;
        RECT 53.520 -1.345 53.690 0.000 ;
        RECT 54.400 -1.205 54.570 0.000 ;
        RECT 54.750 -0.215 55.080 0.000 ;
        RECT 55.280 -1.345 55.450 0.000 ;
        RECT 55.830 -1.345 56.000 0.000 ;
        RECT 56.710 -1.205 56.880 0.000 ;
        RECT 57.590 -1.345 57.760 0.000 ;
        RECT 58.470 -1.205 58.640 0.000 ;
        RECT 59.020 -1.345 59.190 0.000 ;
        RECT 59.900 -1.205 60.070 0.000 ;
        RECT 60.780 -1.345 60.950 0.000 ;
        RECT 68.290 -0.095 70.005 0.000 ;
        RECT 72.315 -0.095 74.335 0.000 ;
        RECT 66.380 -0.575 67.270 -0.405 ;
        RECT 67.550 -0.575 68.220 -0.405 ;
        RECT 66.380 -0.795 66.910 -0.785 ;
        RECT 66.380 -0.955 66.965 -0.795 ;
        RECT 1.485 -1.500 1.655 -1.390 ;
        RECT 2.550 -1.705 60.990 -1.535 ;
        RECT 64.375 -1.785 66.075 -1.035 ;
        RECT 66.795 -1.805 66.965 -0.955 ;
        RECT 67.325 -1.805 67.495 -0.795 ;
        RECT 67.855 -0.815 68.025 -0.795 ;
        RECT 67.855 -0.985 68.385 -0.815 ;
        RECT 67.855 -1.805 68.025 -0.985 ;
      LAYER met1 ;
        RECT 0.000 178.940 80.000 197.965 ;
        RECT 0.000 176.865 80.020 178.940 ;
        RECT 0.000 168.055 80.000 176.865 ;
        RECT -0.115 129.240 80.145 168.055 ;
        RECT 0.000 128.185 80.000 129.240 ;
        RECT -0.115 93.860 80.145 128.185 ;
        RECT 0.000 92.545 80.000 93.860 ;
        RECT 0.000 89.445 80.060 92.545 ;
        RECT -0.145 87.715 80.060 89.445 ;
        RECT 0.000 78.600 80.060 87.715 ;
        RECT -0.115 70.895 80.060 78.600 ;
        POLYGON 80.060 70.950 80.115 70.895 80.060 70.895 ;
        RECT -0.115 55.155 80.115 70.895 ;
        RECT 0.000 49.185 80.115 55.155 ;
        RECT 0.000 33.690 80.000 49.185 ;
        RECT 0.000 28.085 80.115 33.690 ;
        RECT 0.000 22.980 80.000 28.085 ;
        RECT 0.000 17.450 80.115 22.980 ;
        RECT 0.000 0.000 80.000 17.450 ;
        RECT 0.260 -0.130 0.520 0.000 ;
        POLYGON 1.045 -0.100 1.045 -0.130 1.015 -0.130 ;
        RECT 1.045 -0.130 1.275 0.000 ;
        POLYGON 1.015 -0.130 1.015 -0.240 0.905 -0.240 ;
        RECT 1.015 -0.200 1.275 -0.130 ;
        RECT 1.015 -0.240 1.235 -0.200 ;
        POLYGON 1.235 -0.200 1.275 -0.200 1.235 -0.240 ;
        POLYGON 0.905 -0.240 0.905 -0.470 0.675 -0.470 ;
        RECT 0.675 -1.465 0.905 -0.470 ;
        POLYGON 0.905 -0.240 1.235 -0.240 0.905 -0.570 ;
        RECT 1.460 -0.610 1.690 0.000 ;
        POLYGON 1.690 -0.235 2.065 -0.610 1.690 -0.610 ;
        RECT 2.140 -0.255 2.370 0.000 ;
        RECT 3.880 -0.080 30.555 0.000 ;
        POLYGON 33.830 0.000 33.910 0.000 33.910 -0.080 ;
        RECT 33.910 -0.080 34.315 0.000 ;
        POLYGON 22.755 -0.080 22.760 -0.080 22.760 -0.085 ;
        RECT 22.760 -0.085 23.425 -0.080 ;
        POLYGON 2.370 -0.085 2.540 -0.255 2.370 -0.255 ;
        POLYGON 22.760 -0.085 22.785 -0.085 22.785 -0.110 ;
        RECT 22.785 -0.110 23.425 -0.085 ;
        POLYGON 23.425 -0.080 23.455 -0.080 23.425 -0.110 ;
        POLYGON 33.910 -0.080 33.940 -0.080 33.940 -0.110 ;
        RECT 33.940 -0.110 34.315 -0.080 ;
        POLYGON 35.570 0.000 35.655 0.000 35.655 -0.085 ;
        RECT 35.655 -0.085 42.895 0.000 ;
        POLYGON 42.895 0.000 42.980 0.000 42.895 -0.085 ;
        POLYGON 43.390 0.000 43.390 -0.085 43.305 -0.085 ;
        RECT 43.390 -0.085 47.720 0.000 ;
        POLYGON 33.940 -0.110 34.085 -0.110 34.085 -0.255 ;
        RECT 2.140 -0.485 18.040 -0.255 ;
        POLYGON 17.370 -0.485 17.400 -0.485 17.400 -0.515 ;
        RECT 17.400 -0.515 18.040 -0.485 ;
        RECT 21.550 -0.540 29.630 -0.280 ;
        RECT 29.770 -0.535 32.915 -0.275 ;
        RECT 34.085 -0.325 34.315 -0.110 ;
        POLYGON 43.305 -0.085 43.305 -0.225 43.165 -0.225 ;
        RECT 43.305 -0.190 47.720 -0.085 ;
        RECT 43.305 -0.225 43.370 -0.190 ;
        RECT 35.460 -0.485 38.120 -0.225 ;
        POLYGON 43.165 -0.225 43.165 -0.350 43.040 -0.350 ;
        RECT 43.165 -0.350 43.370 -0.225 ;
        POLYGON 43.370 -0.190 43.530 -0.190 43.370 -0.350 ;
        POLYGON 47.580 -0.190 47.680 -0.190 47.680 -0.290 ;
        RECT 47.680 -0.290 47.720 -0.190 ;
        POLYGON 47.720 0.000 48.010 -0.290 47.720 -0.290 ;
        POLYGON 54.810 -0.120 54.810 -0.290 54.640 -0.290 ;
        RECT 54.810 -0.290 55.040 0.000 ;
        RECT 56.680 -0.145 56.910 0.000 ;
        POLYGON 47.680 -0.290 47.740 -0.290 47.740 -0.350 ;
        RECT 47.740 -0.350 55.040 -0.290 ;
        RECT 39.390 -0.610 43.110 -0.350 ;
        POLYGON 43.110 -0.350 43.370 -0.350 43.110 -0.610 ;
        RECT 45.040 -0.610 47.515 -0.350 ;
        POLYGON 47.740 -0.350 47.910 -0.350 47.910 -0.520 ;
        RECT 47.910 -0.520 55.040 -0.350 ;
        RECT 1.460 -0.750 2.065 -0.610 ;
        POLYGON 2.065 -0.610 2.205 -0.750 2.065 -0.750 ;
        RECT 62.430 -0.730 62.690 -0.120 ;
        RECT 63.680 -0.595 64.880 0.000 ;
        POLYGON 65.530 0.000 65.635 0.000 65.635 -0.105 ;
        RECT 1.460 -1.765 61.195 -0.750 ;
        RECT 65.635 -0.845 65.775 0.000 ;
        POLYGON 66.830 -0.080 66.830 -0.375 66.535 -0.375 ;
        RECT 66.830 -0.375 67.095 0.000 ;
        RECT 66.320 -0.605 67.095 -0.375 ;
        RECT 67.355 -0.375 67.495 0.000 ;
        POLYGON 68.000 0.000 68.080 0.000 68.080 -0.080 ;
        RECT 68.080 -0.080 68.215 0.000 ;
        POLYGON 68.215 0.000 68.295 -0.080 68.215 -0.080 ;
        POLYGON 68.080 -0.080 68.215 -0.080 68.215 -0.215 ;
        RECT 68.215 -0.215 68.295 -0.080 ;
        POLYGON 67.495 -0.215 67.655 -0.375 67.495 -0.375 ;
        POLYGON 68.215 -0.215 68.295 -0.215 68.295 -0.295 ;
        POLYGON 68.295 -0.080 68.510 -0.295 68.295 -0.295 ;
        POLYGON 68.295 -0.295 68.370 -0.295 68.370 -0.370 ;
        RECT 67.355 -0.605 68.155 -0.375 ;
        POLYGON 68.370 -0.605 68.370 -0.705 68.270 -0.705 ;
        RECT 68.370 -0.705 68.510 -0.295 ;
        POLYGON 65.775 -0.705 65.915 -0.845 65.775 -0.845 ;
        POLYGON 68.270 -0.705 68.270 -0.755 68.220 -0.755 ;
        RECT 68.270 -0.755 68.510 -0.705 ;
        POLYGON 66.320 -0.755 66.320 -0.845 66.230 -0.845 ;
        RECT 66.320 -0.845 66.970 -0.755 ;
        POLYGON 68.220 -0.755 68.220 -0.785 68.190 -0.785 ;
        RECT 68.220 -0.785 68.510 -0.755 ;
        RECT 65.635 -0.985 66.970 -0.845 ;
        RECT 67.795 -1.015 68.510 -0.785 ;
        POLYGON 79.110 -0.915 79.110 -1.015 79.010 -1.015 ;
        RECT 79.110 -1.015 79.370 -0.835 ;
        POLYGON 79.010 -1.015 79.010 -1.125 78.900 -1.125 ;
        RECT 79.010 -1.125 79.370 -1.015 ;
        RECT 64.375 -1.775 67.525 -1.125 ;
        POLYGON 78.900 -1.125 78.900 -1.195 78.830 -1.195 ;
        RECT 78.900 -1.195 79.370 -1.125 ;
        RECT 75.255 -1.475 79.370 -1.195 ;
      LAYER met2 ;
        RECT 0.210 176.115 79.915 197.965 ;
        RECT 0.210 4.670 79.435 176.115 ;
        RECT 0.210 3.595 22.075 4.670 ;
        RECT 0.210 2.720 12.475 3.595 ;
        RECT 0.210 0.000 3.095 2.720 ;
        RECT 3.885 0.000 5.140 2.720 ;
        RECT 5.930 0.000 12.475 2.720 ;
        RECT 13.295 0.565 22.075 3.595 ;
        RECT 13.295 0.000 16.030 0.565 ;
        RECT 16.850 0.000 22.075 0.565 ;
        RECT 22.895 3.335 79.435 4.670 ;
        RECT 22.895 2.315 44.965 3.335 ;
        RECT 22.895 0.950 28.210 2.315 ;
        RECT 22.895 0.150 26.320 0.950 ;
        RECT 22.785 0.000 26.320 0.150 ;
        RECT 27.140 0.000 28.210 0.950 ;
        RECT 29.030 1.585 44.965 2.315 ;
        RECT 29.030 0.510 31.535 1.585 ;
        RECT 29.030 0.000 30.470 0.510 ;
        RECT 31.290 0.000 31.535 0.510 ;
        RECT 32.355 1.335 44.965 1.585 ;
        RECT 32.355 0.720 38.110 1.335 ;
        RECT 32.355 0.000 38.120 0.720 ;
        RECT 38.930 0.000 44.965 1.335 ;
        RECT 45.785 0.515 79.435 3.335 ;
        RECT 45.785 0.000 67.995 0.515 ;
        RECT 69.205 0.300 79.435 0.515 ;
        RECT 69.205 0.000 76.000 0.300 ;
        RECT 77.200 0.020 79.435 0.300 ;
        RECT 76.920 0.000 79.435 0.020 ;
        RECT 0.260 -1.065 0.520 0.000 ;
        RECT 1.080 -0.340 1.380 0.000 ;
        POLYGON 1.380 0.000 1.720 -0.340 1.380 -0.340 ;
        POLYGON 0.260 -1.065 0.520 -1.065 0.520 -1.325 ;
        POLYGON 0.520 -0.955 0.680 -1.115 0.520 -1.115 ;
        RECT 1.080 -1.110 1.720 -0.340 ;
        RECT 0.520 -1.325 0.680 -1.115 ;
        POLYGON 0.520 -1.325 0.670 -1.325 0.670 -1.475 ;
        RECT 0.670 -1.475 0.680 -1.325 ;
        POLYGON 0.680 -1.115 1.040 -1.475 0.680 -1.475 ;
        POLYGON 0.670 -1.475 0.930 -1.475 0.930 -1.735 ;
        RECT 0.930 -1.735 2.160 -1.475 ;
        RECT 2.365 -1.735 3.005 0.000 ;
        POLYGON 6.615 0.000 6.615 -0.020 6.595 -0.020 ;
        RECT 6.615 -0.020 6.965 0.000 ;
        POLYGON 6.965 0.000 6.985 0.000 6.965 -0.020 ;
        POLYGON 6.595 -0.020 6.595 -0.390 6.225 -0.390 ;
        POLYGON 6.595 -0.020 6.965 -0.020 6.595 -0.390 ;
        POLYGON 17.600 -0.080 17.600 -0.255 17.425 -0.255 ;
        RECT 17.600 -0.255 17.860 0.000 ;
        POLYGON 17.860 -0.080 18.035 -0.255 17.860 -0.255 ;
        POLYGON 6.225 -0.390 6.225 -0.485 6.130 -0.485 ;
        RECT 6.225 -0.485 6.500 -0.390 ;
        POLYGON 6.500 -0.390 6.595 -0.390 6.500 -0.485 ;
        POLYGON 6.390 -0.485 6.500 -0.485 6.390 -0.595 ;
        RECT 17.400 -0.515 18.040 -0.255 ;
        RECT 6.895 -1.765 10.715 -0.755 ;
        RECT 19.235 -1.765 21.375 0.000 ;
        POLYGON 21.775 -0.110 21.775 -0.280 21.605 -0.280 ;
        RECT 21.775 -0.280 22.035 0.000 ;
        RECT 22.785 -0.110 23.425 0.000 ;
        POLYGON 24.045 0.000 24.045 -0.110 23.935 -0.110 ;
        RECT 24.045 -0.110 26.265 0.000 ;
        POLYGON 23.935 -0.110 23.935 -0.125 23.920 -0.125 ;
        RECT 23.935 -0.125 26.265 -0.110 ;
        POLYGON 22.035 -0.125 22.190 -0.280 22.035 -0.280 ;
        POLYGON 23.920 -0.125 23.920 -0.150 23.895 -0.150 ;
        RECT 23.920 -0.150 26.265 -0.125 ;
        RECT 21.550 -0.540 22.190 -0.280 ;
        POLYGON 23.895 -0.150 23.895 -0.350 23.695 -0.350 ;
        RECT 23.895 -0.350 26.265 -0.150 ;
        POLYGON 23.695 -0.350 23.695 -0.540 23.505 -0.540 ;
        RECT 23.695 -0.540 26.265 -0.350 ;
        POLYGON 29.085 -0.185 29.085 -0.280 28.990 -0.280 ;
        RECT 29.085 -0.280 29.350 0.000 ;
        POLYGON 29.350 0.000 29.630 -0.280 29.350 -0.280 ;
        RECT 28.990 -0.540 29.630 -0.280 ;
        RECT 29.770 -0.535 30.410 0.000 ;
        POLYGON 32.355 -0.085 32.355 -0.165 32.275 -0.165 ;
        RECT 32.355 -0.165 32.615 0.000 ;
        RECT 32.275 -0.275 32.615 -0.165 ;
        POLYGON 32.615 -0.085 32.805 -0.275 32.615 -0.275 ;
        RECT 32.275 -0.535 32.915 -0.275 ;
        POLYGON 23.505 -0.540 23.505 -0.750 23.295 -0.750 ;
        RECT 23.505 -0.750 26.265 -0.540 ;
        RECT 22.995 -1.760 26.265 -0.750 ;
        RECT 33.400 -1.765 34.670 0.000 ;
        POLYGON 35.325 0.000 35.350 0.000 35.350 -0.025 ;
        RECT 35.350 -0.025 35.695 0.000 ;
        POLYGON 35.695 0.000 35.720 -0.025 35.695 -0.025 ;
        POLYGON 37.705 0.000 37.705 -0.025 37.680 -0.025 ;
        RECT 37.705 -0.025 38.120 0.000 ;
        POLYGON 35.350 -0.025 35.460 -0.025 35.460 -0.135 ;
        RECT 35.460 -0.225 35.720 -0.025 ;
        POLYGON 35.720 -0.025 35.920 -0.225 35.720 -0.225 ;
        POLYGON 37.680 -0.025 37.680 -0.225 37.480 -0.225 ;
        RECT 37.680 -0.225 38.120 -0.025 ;
        RECT 35.460 -0.485 36.100 -0.225 ;
        RECT 37.480 -0.485 38.120 -0.225 ;
        POLYGON 39.770 -0.005 39.770 -0.350 39.425 -0.350 ;
        RECT 39.770 -0.350 40.030 0.000 ;
        POLYGON 42.060 0.000 42.060 -0.310 41.750 -0.310 ;
        RECT 42.060 -0.310 42.120 0.000 ;
        POLYGON 42.120 0.000 42.430 0.000 42.120 -0.310 ;
        POLYGON 47.375 -0.180 47.375 -0.310 47.245 -0.310 ;
        RECT 47.375 -0.310 47.515 0.000 ;
        RECT 49.395 -0.165 50.165 0.000 ;
        POLYGON 35.720 -0.485 35.920 -0.485 35.720 -0.685 ;
        RECT 39.390 -0.610 40.030 -0.350 ;
        POLYGON 41.750 -0.310 41.750 -0.610 41.450 -0.610 ;
        POLYGON 41.450 -0.610 41.450 -0.680 41.380 -0.680 ;
        RECT 41.450 -0.680 41.750 -0.610 ;
        POLYGON 41.750 -0.310 42.120 -0.310 41.750 -0.680 ;
        POLYGON 47.245 -0.310 47.245 -0.350 47.205 -0.350 ;
        RECT 47.245 -0.350 47.515 -0.310 ;
        RECT 46.770 -0.610 47.515 -0.350 ;
        POLYGON 51.970 -0.330 51.970 -0.570 51.730 -0.570 ;
        RECT 51.970 -0.570 52.230 0.000 ;
        RECT 52.525 -0.040 54.155 0.000 ;
        POLYGON 52.525 -0.040 52.825 -0.040 52.825 -0.340 ;
        RECT 52.825 -0.340 54.155 -0.040 ;
        POLYGON 52.230 -0.340 52.460 -0.570 52.230 -0.570 ;
        POLYGON 41.380 -0.680 41.380 -0.685 41.375 -0.685 ;
        RECT 41.380 -0.685 41.530 -0.680 ;
        POLYGON 41.375 -0.685 41.375 -0.705 41.355 -0.705 ;
        RECT 41.375 -0.705 41.530 -0.685 ;
        POLYGON 38.650 -0.705 38.845 -0.900 38.650 -0.900 ;
        POLYGON 41.355 -0.705 41.355 -0.900 41.160 -0.900 ;
        RECT 41.355 -0.900 41.530 -0.705 ;
        POLYGON 41.530 -0.680 41.750 -0.680 41.530 -0.900 ;
        RECT 51.690 -0.850 52.460 -0.570 ;
        POLYGON 52.825 -0.340 53.335 -0.340 53.335 -0.850 ;
        RECT 53.335 -0.850 54.155 -0.340 ;
        POLYGON 53.335 -0.850 53.385 -0.850 53.385 -0.900 ;
        RECT 53.385 -0.900 54.155 -0.850 ;
        RECT 38.650 -1.160 41.270 -0.900 ;
        POLYGON 41.270 -0.900 41.530 -0.900 41.270 -1.160 ;
        POLYGON 53.385 -0.900 53.645 -0.900 53.645 -1.160 ;
        RECT 53.645 -0.985 54.155 -0.900 ;
        POLYGON 54.155 -0.185 54.955 -0.985 54.155 -0.985 ;
        RECT 62.430 -0.760 62.690 0.000 ;
        RECT 63.680 -0.595 64.385 0.000 ;
        POLYGON 76.920 0.000 77.330 0.000 76.920 -0.410 ;
        RECT 66.540 -0.840 67.360 -0.560 ;
        POLYGON 66.540 -0.840 66.685 -0.840 66.685 -0.985 ;
        RECT 66.685 -0.985 66.835 -0.840 ;
        RECT 53.645 -1.160 65.200 -0.985 ;
        POLYGON 66.685 -0.985 66.835 -0.985 66.835 -1.135 ;
        POLYGON 67.095 -0.840 67.360 -0.840 67.095 -1.105 ;
        RECT 77.390 -0.850 78.210 -0.570 ;
        POLYGON 78.710 -0.815 78.710 -0.820 78.705 -0.820 ;
        RECT 78.710 -0.820 78.910 0.000 ;
        POLYGON 77.410 -0.850 77.610 -0.850 77.610 -1.050 ;
        RECT 77.870 -1.050 77.980 -0.850 ;
        POLYGON 77.980 -0.850 78.180 -0.850 77.980 -1.050 ;
        RECT 78.905 -0.905 78.910 -0.820 ;
        POLYGON 78.905 -0.905 78.910 -0.905 78.905 -0.910 ;
        RECT 77.870 -1.105 77.925 -1.050 ;
        POLYGON 77.925 -1.050 77.980 -1.050 77.925 -1.105 ;
        RECT 77.870 -1.135 77.895 -1.105 ;
        POLYGON 77.895 -1.105 77.925 -1.105 77.895 -1.135 ;
        POLYGON 77.870 -1.135 77.895 -1.135 77.870 -1.160 ;
        POLYGON 38.650 -1.160 38.845 -1.160 38.650 -1.355 ;
        POLYGON 53.645 -1.160 53.695 -1.160 53.695 -1.210 ;
        RECT 53.695 -1.210 65.200 -1.160 ;
        RECT 49.590 -1.490 50.360 -1.210 ;
        POLYGON 49.590 -1.490 49.855 -1.490 49.855 -1.755 ;
        POLYGON 50.115 -1.490 50.360 -1.490 50.115 -1.735 ;
        POLYGON 53.695 -1.210 54.155 -1.210 54.155 -1.670 ;
        RECT 54.155 -1.670 65.200 -1.210 ;
        RECT 75.125 -1.475 75.895 -1.195 ;
        RECT 79.110 -1.475 79.370 0.000 ;
        POLYGON 54.155 -1.670 54.220 -1.670 54.220 -1.735 ;
        RECT 54.220 -1.735 65.200 -1.670 ;
        POLYGON 54.220 -1.735 54.240 -1.735 54.240 -1.755 ;
        RECT 54.240 -1.755 65.200 -1.735 ;
        POLYGON 54.240 -1.755 54.250 -1.755 54.250 -1.765 ;
        RECT 54.250 -1.765 65.200 -1.755 ;
        POLYGON 54.250 -1.765 54.270 -1.765 54.270 -1.785 ;
        RECT 54.270 -1.785 65.200 -1.765 ;
      LAYER met3 ;
        RECT 0.400 187.925 79.570 197.965 ;
        RECT 0.400 183.140 78.840 187.925 ;
        RECT 0.400 176.850 78.180 183.140 ;
        RECT 1.420 35.170 78.180 176.850 ;
        RECT 1.420 0.000 45.465 35.170 ;
        RECT 46.595 8.070 78.180 35.170 ;
        RECT 46.595 0.000 62.420 8.070 ;
        RECT 64.290 0.000 78.180 8.070 ;
        RECT 1.415 -1.090 2.205 -0.360 ;
        POLYGON 3.680 -1.125 3.680 -1.175 3.630 -1.175 ;
        RECT 3.680 -1.175 4.010 0.000 ;
        POLYGON 4.010 -0.775 4.410 -1.175 4.010 -1.175 ;
        RECT 3.630 -1.495 4.410 -1.175 ;
        RECT 6.455 -1.790 10.715 0.000 ;
        RECT 22.635 -1.785 27.635 0.000 ;
        RECT 49.415 -0.190 53.035 0.000 ;
        POLYGON 53.035 0.000 53.225 -0.190 53.035 -0.190 ;
        POLYGON 52.755 -0.190 53.110 -0.190 53.110 -0.545 ;
        RECT 53.110 -0.545 53.225 -0.190 ;
        POLYGON 53.225 -0.190 53.580 -0.545 53.225 -0.545 ;
        POLYGON 65.510 -0.310 65.510 -0.545 65.275 -0.545 ;
        RECT 65.510 -0.545 65.815 0.000 ;
        POLYGON 77.075 0.000 77.075 -0.415 76.660 -0.415 ;
        RECT 77.075 -0.415 77.110 0.000 ;
        POLYGON 77.110 0.000 77.525 0.000 77.110 -0.415 ;
        POLYGON 76.660 -0.415 76.660 -0.535 76.540 -0.535 ;
        RECT 51.685 -0.875 52.465 -0.545 ;
        POLYGON 53.110 -0.545 53.225 -0.545 53.225 -0.660 ;
        RECT 53.225 -0.660 54.320 -0.545 ;
        POLYGON 53.225 -0.660 53.430 -0.660 53.430 -0.865 ;
        RECT 53.430 -0.865 54.320 -0.660 ;
        POLYGON 55.510 -0.545 55.510 -0.865 55.190 -0.865 ;
        RECT 55.510 -0.865 56.785 -0.545 ;
        RECT 65.035 -0.865 65.815 -0.545 ;
        RECT 66.560 -0.865 67.340 -0.535 ;
        POLYGON 76.540 -0.535 76.540 -0.545 76.530 -0.545 ;
        RECT 76.540 -0.545 76.660 -0.535 ;
        RECT 75.120 -0.865 76.660 -0.545 ;
        POLYGON 76.660 -0.415 77.110 -0.415 76.660 -0.865 ;
        POLYGON 55.190 -0.865 55.190 -0.875 55.180 -0.875 ;
        RECT 55.190 -0.875 55.510 -0.865 ;
        POLYGON 55.180 -0.875 55.180 -0.995 55.060 -0.995 ;
        RECT 55.180 -0.995 55.510 -0.875 ;
        POLYGON 55.510 -0.865 55.640 -0.865 55.510 -0.995 ;
        RECT 77.410 -0.875 78.190 -0.545 ;
        POLYGON 55.060 -0.995 55.060 -1.185 54.870 -1.185 ;
        RECT 55.060 -1.185 55.205 -0.995 ;
        RECT 49.610 -1.300 55.205 -1.185 ;
        POLYGON 55.205 -0.995 55.510 -0.995 55.205 -1.300 ;
        RECT 49.610 -1.505 55.000 -1.300 ;
        POLYGON 55.000 -1.300 55.205 -1.300 55.000 -1.505 ;
        RECT 75.145 -1.500 75.925 -1.170 ;
        RECT 49.610 -1.515 50.340 -1.505 ;
        POLYGON 50.340 -1.505 50.350 -1.505 50.340 -1.515 ;
      LAYER met4 ;
        RECT 1.670 173.350 78.330 197.965 ;
        RECT 0.965 93.365 78.970 173.350 ;
        RECT 1.670 67.600 78.330 93.365 ;
        RECT 0.965 66.900 78.970 67.600 ;
        RECT 1.670 61.650 78.330 66.900 ;
        RECT 0.965 61.050 78.970 61.650 ;
        RECT 1.670 55.800 78.330 61.050 ;
        RECT 0.965 55.100 78.970 55.800 ;
        RECT 3.010 54.470 46.690 55.100 ;
        RECT 36.840 50.690 38.360 54.470 ;
        RECT 1.670 49.710 78.330 50.690 ;
        RECT 52.545 46.430 54.065 49.710 ;
        RECT 3.010 45.300 46.690 45.930 ;
        RECT 0.965 44.600 78.970 45.300 ;
        RECT 1.670 39.150 78.330 44.600 ;
        RECT 0.965 38.550 78.970 39.150 ;
        RECT 1.670 34.300 78.330 38.550 ;
        RECT 0.965 33.700 78.970 34.300 ;
        RECT 1.670 29.450 78.330 33.700 ;
        RECT 0.965 28.850 78.970 29.450 ;
        RECT 1.670 23.400 78.330 28.850 ;
        RECT 0.965 22.800 78.970 23.400 ;
        RECT 1.670 17.350 78.330 22.800 ;
        RECT 0.965 16.750 78.970 17.350 ;
        RECT 1.365 12.500 78.570 16.750 ;
        RECT 0.965 11.900 78.970 12.500 ;
        RECT 1.670 6.450 78.330 11.900 ;
        RECT 0.965 5.850 78.970 6.450 ;
        RECT 1.670 0.000 78.330 5.850 ;
        RECT 1.450 -0.870 52.440 -0.540 ;
        RECT 53.565 -0.870 56.760 -0.540 ;
        RECT 65.060 -0.870 67.315 -0.540 ;
        RECT 75.145 -0.870 78.165 -0.540 ;
        RECT 3.655 -1.500 75.900 -1.170 ;
      LAYER met5 ;
        RECT 0.000 166.575 80.000 197.965 ;
        RECT 0.000 100.925 9.600 166.575 ;
        RECT 75.400 100.925 80.000 166.575 ;
        RECT 0.000 94.550 80.000 100.925 ;
        RECT 2.870 16.250 77.130 94.550 ;
        RECT 2.565 13.000 77.370 16.250 ;
        RECT 2.870 0.100 77.130 13.000 ;
  END
END sky130_ef_io__gpiov2_pad
END LIBRARY

