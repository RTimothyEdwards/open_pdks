magic
tech sky130A
magscale 1 2
timestamp 1607710972
<< metal1 >>
rect 15049 7630 17239 7665
rect 15049 6925 15080 7630
rect 17210 6925 17239 7630
rect 15049 6891 17239 6925
rect 4185 -163 10707 -7
rect 15240 -163 17187 6891
rect 4185 -1307 17187 -163
rect 4185 -2107 16387 -1307
tri 16387 -2107 17187 -1307 nw
<< via1 >>
rect 15080 6925 17210 7630
<< metal2 >>
rect 132 38667 2749 38676
rect 132 34800 141 38667
rect 2740 34800 2749 38667
rect 132 34791 2749 34800
rect 14940 8809 17228 8840
rect 14940 7939 15154 8809
rect 16192 7939 17228 8809
rect 14940 7910 17228 7939
rect 15049 7630 17239 7665
rect 15049 6925 15080 7630
rect 17210 7605 17239 7630
rect 17213 6966 17239 7605
rect 17210 6925 17239 6966
rect 15049 6891 17239 6925
<< via2 >>
rect 141 34800 2740 38667
rect 15154 7939 16192 8809
rect 15116 6966 17210 7605
rect 17210 6966 17213 7605
<< metal3 >>
rect 102 38667 2772 38714
rect 102 34800 141 38667
rect 2740 34800 2772 38667
rect 102 34753 2772 34800
rect 15121 8809 17228 8840
rect 15121 7939 15154 8809
rect 17192 7939 17228 8809
rect 15121 7910 17228 7939
rect 15088 7605 17228 7632
rect 15088 6966 15116 7605
rect 17213 6966 17228 7605
rect 15088 6939 17228 6966
rect 5228 2263 7341 2269
rect 5228 1400 5234 2263
rect 7335 1400 7341 2263
rect 5228 1394 7341 1400
rect 7705 2261 9818 2267
rect 7705 1398 7711 2261
rect 9812 1398 9818 2261
rect 7705 1392 9818 1398
<< via3 >>
rect 141 34800 2740 38667
rect 15154 7939 16192 8809
rect 16192 7939 17192 8809
rect 15116 6966 17213 7605
rect 5234 1400 7335 2263
rect 7711 1398 9812 2261
<< metal4 >>
rect 132 38667 2749 38676
rect 132 34800 141 38667
rect 2740 34800 2749 38667
rect 132 34791 2749 34800
rect 14940 8809 17228 8840
rect 14940 7939 15154 8809
rect 17192 7939 17228 8809
rect 14940 7910 17228 7939
rect 14985 7605 17233 7630
rect 14985 6966 15116 7605
rect 17213 6966 17233 7605
rect 14985 6940 17233 6966
rect 5228 2263 7341 2269
rect 5228 1400 5234 2263
rect 7335 1400 7341 2263
rect 5228 1394 7341 1400
rect 7705 2261 9818 2267
rect 7705 1398 7711 2261
rect 9812 1398 9818 2261
rect 7705 1392 9818 1398
<< properties >>
string FIXED_BBOX 0 -7 15000 39593
<< end >>
