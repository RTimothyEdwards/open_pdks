magic
tech sky130A
magscale 1 2
timestamp 1602597384
<< error_s >>
rect 14469 39226 14535 39242
rect 3098 36629 3170 38629
rect 3369 36662 3487 38556
rect 3758 36629 3818 38629
rect 4018 36629 4090 38629
rect 4289 36662 4407 38556
rect 4678 36629 4738 38629
rect 4938 36629 5010 38629
rect 5209 36662 5327 38556
rect 5598 36629 5658 38629
rect 5858 36629 5930 38629
rect 6129 36662 6247 38556
rect 6518 36629 6578 38629
rect 6778 36629 6850 38629
rect 7049 36662 7167 38556
rect 7438 36629 7498 38629
rect 7698 36629 7770 38629
rect 7969 36662 8087 38556
rect 8358 36629 8418 38629
rect 8618 36629 8690 38629
rect 8889 36662 9007 38556
rect 9278 36629 9338 38629
rect 9538 36629 9610 38629
rect 9809 36662 9927 38556
rect 10198 36629 10258 38629
rect 10458 36629 10530 38629
rect 10729 36662 10847 38556
rect 11118 36629 11178 38629
rect 11378 36629 11450 38629
rect 11649 36662 11767 38556
rect 12038 36629 12098 38629
rect 12298 36629 12370 38629
rect 12569 36662 12687 38556
rect 12958 36629 13018 38629
rect 3098 32029 3170 36029
rect 3369 32062 3487 35996
rect 3758 32029 3818 36029
rect 4018 32029 4090 36029
rect 4289 32062 4407 35996
rect 4678 32029 4738 36029
rect 4938 32029 5010 36029
rect 5209 32062 5327 35996
rect 5598 32029 5658 36029
rect 5858 32029 5930 36029
rect 6129 32062 6247 35996
rect 6518 32029 6578 36029
rect 6778 32029 6850 36029
rect 7049 32062 7167 35996
rect 7438 32029 7498 36029
rect 7698 32029 7770 36029
rect 7969 32062 8087 35996
rect 8358 32029 8418 36029
rect 8618 32029 8690 36029
rect 8889 32062 9007 35996
rect 9278 32029 9338 36029
rect 9538 32029 9610 36029
rect 9809 32062 9927 35996
rect 10198 32029 10258 36029
rect 10458 32029 10530 36029
rect 10729 32062 10847 35996
rect 11118 32029 11178 36029
rect 11378 32029 11450 36029
rect 11649 32062 11767 35996
rect 12038 32029 12098 36029
rect 12298 32029 12370 36029
rect 12569 32062 12687 35996
rect 12958 32029 13018 36029
rect 3098 27429 3170 31429
rect 3369 27462 3487 31396
rect 3758 27429 3818 31429
rect 4018 27429 4090 31429
rect 4289 27462 4407 31396
rect 4678 27429 4738 31429
rect 4938 27429 5010 31429
rect 5209 27462 5327 31396
rect 5598 27429 5658 31429
rect 5858 27429 5930 31429
rect 6129 27462 6247 31396
rect 6518 27429 6578 31429
rect 6778 27429 6850 31429
rect 7049 27462 7167 31396
rect 7438 27429 7498 31429
rect 7698 27429 7770 31429
rect 7969 27462 8087 31396
rect 8358 27429 8418 31429
rect 8618 27429 8690 31429
rect 8889 27462 9007 31396
rect 9278 27429 9338 31429
rect 9538 27429 9610 31429
rect 9809 27462 9927 31396
rect 10198 27429 10258 31429
rect 10458 27429 10530 31429
rect 10729 27462 10847 31396
rect 11118 27429 11178 31429
rect 11378 27429 11450 31429
rect 11649 27462 11767 31396
rect 12038 27429 12098 31429
rect 12298 27429 12370 31429
rect 12569 27462 12687 31396
rect 12958 27429 13018 31429
rect 4938 22829 5010 26829
rect 5209 22862 5327 26796
rect 5598 22829 5658 26829
rect 5858 22829 5930 26829
rect 6129 22862 6247 26796
rect 6518 22829 6578 26829
rect 6778 22829 6850 26829
rect 7049 22862 7167 26796
rect 7438 22829 7498 26829
rect 7698 22829 7770 26829
rect 7969 22862 8087 26796
rect 8358 22829 8418 26829
rect 8618 22829 8690 26829
rect 8889 22862 9007 26796
rect 9278 22829 9338 26829
rect 9538 22829 9610 26829
rect 9809 22862 9927 26796
rect 10198 22829 10258 26829
rect 10458 22829 10530 26829
rect 10729 22862 10847 26796
rect 11118 22829 11178 26829
rect 11378 22829 11450 26829
rect 11649 22862 11767 26796
rect 12038 22829 12098 26829
rect 12298 22829 12370 26829
rect 12569 22862 12687 26796
rect 12958 22829 13018 26829
rect 4938 18229 5010 22229
rect 5209 18262 5327 22196
rect 5598 18229 5658 22229
rect 5858 18229 5930 22229
rect 6129 18262 6247 22196
rect 6518 18229 6578 22229
rect 6778 18229 6850 22229
rect 7049 18262 7167 22196
rect 7438 18229 7498 22229
rect 7698 18229 7770 22229
rect 7969 18262 8087 22196
rect 8358 18229 8418 22229
rect 8618 18229 8690 22229
rect 8889 18262 9007 22196
rect 9278 18229 9338 22229
rect 9538 18229 9610 22229
rect 9809 18262 9927 22196
rect 10198 18229 10258 22229
rect 10458 18229 10530 22229
rect 10729 18262 10847 22196
rect 11118 18229 11178 22229
rect 11378 18229 11450 22229
rect 11649 18262 11767 22196
rect 12038 18229 12098 22229
rect 12298 18229 12370 22229
rect 12569 18262 12687 22196
rect 12958 18229 13018 22229
rect 1900 14464 1966 14480
rect 3682 14470 3748 14486
rect 4938 13629 5010 17629
rect 5209 13662 5327 17596
rect 5598 13629 5658 17629
rect 5858 13629 5930 17629
rect 6129 13662 6247 17596
rect 6518 13629 6578 17629
rect 6778 13629 6850 17629
rect 7049 13662 7167 17596
rect 7438 13629 7498 17629
rect 7698 13629 7770 17629
rect 7969 13662 8087 17596
rect 8358 13629 8418 17629
rect 8618 13629 8690 17629
rect 8889 13662 9007 17596
rect 9278 13629 9338 17629
rect 9538 13629 9610 17629
rect 9809 13662 9927 17596
rect 10198 13629 10258 17629
rect 10458 13629 10530 17629
rect 10729 13662 10847 17596
rect 11118 13629 11178 17629
rect 11378 13629 11450 17629
rect 11649 13662 11767 17596
rect 12038 13629 12098 17629
rect 12298 13629 12370 17629
rect 12569 13662 12687 17596
rect 12958 13629 13018 17629
rect 3098 9029 3170 13029
rect 3369 9062 3487 12996
rect 3758 9029 3818 13029
rect 4018 9029 4090 13029
rect 4289 9062 4407 12996
rect 4678 9029 4738 13029
rect 4938 9029 5010 13029
rect 5209 9062 5327 12996
rect 5598 9029 5658 13029
rect 5858 9029 5930 13029
rect 6129 9062 6247 12996
rect 6518 9029 6578 13029
rect 6778 9029 6850 13029
rect 7049 9062 7167 12996
rect 7438 9029 7498 13029
rect 7698 9029 7770 13029
rect 7969 9062 8087 12996
rect 8358 9029 8418 13029
rect 8618 9029 8690 13029
rect 8889 9062 9007 12996
rect 9278 9029 9338 13029
rect 9538 9029 9610 13029
rect 9809 9062 9927 12996
rect 10198 9029 10258 13029
rect 10458 9029 10530 13029
rect 10729 9062 10847 12996
rect 11118 9029 11178 13029
rect 11378 9029 11450 13029
rect 11649 9062 11767 12996
rect 12038 9029 12098 13029
rect 12298 9029 12370 13029
rect 12569 9062 12687 12996
rect 12958 9029 13018 13029
rect 214 8281 280 8297
rect 1672 8281 1738 8297
rect 14145 7996 14211 8012
rect 1218 5553 1268 6953
rect 1368 5553 1496 6953
rect 1524 5553 1652 6953
rect 1680 5553 1808 6953
rect 1836 5553 1964 6953
rect 1992 5553 2120 6953
rect 2148 5553 2276 6953
rect 2304 5553 2432 6953
rect 2460 5553 2588 6953
rect 2616 5553 2744 6953
rect 2772 5553 2900 6953
rect 2928 5553 3056 6953
rect 3084 5553 3212 6953
rect 3240 5553 3368 6953
rect 3396 5553 3524 6953
rect 3552 5553 3680 6953
rect 3708 5553 3836 6953
rect 3864 5553 3992 6953
rect 4020 5553 4148 6953
rect 4176 5553 4304 6953
rect 4332 5553 4460 6953
rect 4488 5553 4616 6953
rect 4644 5553 4772 6953
rect 4800 5553 4928 6953
rect 4956 5553 5084 6953
rect 5112 5553 5240 6953
rect 5268 5553 5396 6953
rect 5424 5553 5552 6953
rect 5580 5553 5708 6953
rect 5736 5553 5864 6953
rect 5892 5553 6020 6953
rect 6048 5553 6176 6953
rect 6204 5553 6332 6953
rect 6360 5553 6488 6953
rect 6516 5553 6644 6953
rect 6672 5553 6800 6953
rect 6828 5553 6956 6953
rect 6984 5553 7112 6953
rect 7140 5553 7268 6953
rect 7296 5553 7424 6953
rect 7452 5553 7580 6953
rect 7608 5553 7736 6953
rect 7764 5553 7892 6953
rect 7920 5553 8048 6953
rect 8076 5553 8204 6953
rect 8232 5553 8360 6953
rect 8388 5553 8516 6953
rect 8544 5553 8672 6953
rect 8700 5553 8828 6953
rect 8856 5553 8984 6953
rect 9012 5553 9062 6953
rect 10933 6109 10983 7509
rect 11083 6109 11211 7509
rect 11239 6109 11367 7509
rect 11395 6109 11523 7509
rect 11551 6109 11679 7509
rect 11707 6109 11835 7509
rect 11863 6109 11991 7509
rect 12019 6109 12147 7509
rect 12175 6109 12303 7509
rect 12331 6109 12459 7509
rect 12487 6109 12615 7509
rect 12643 6109 12771 7509
rect 12799 6109 12927 7509
rect 12955 6109 13083 7509
rect 13111 6109 13239 7509
rect 13267 6109 13317 7509
rect 11513 4022 11563 5022
rect 12363 4022 12413 5022
rect 12665 4022 12715 5022
rect 13515 4022 13565 5022
rect 2905 2778 2955 3778
rect 3755 2778 3805 3778
rect 4057 2778 4107 3778
rect 5707 2778 5757 3778
rect 6009 2778 6059 3778
rect 7659 2778 7709 3778
rect 7961 2778 8011 3778
rect 9611 2778 9661 3778
rect 9913 2778 9963 3778
rect 11563 2778 11613 3778
rect 11865 2778 11915 3778
rect 13515 2778 13565 3778
rect 2905 1534 2955 2534
rect 3755 1534 3805 2534
rect 4057 1534 4107 2534
rect 5707 1534 5757 2534
rect 6009 1534 6059 2534
rect 7659 1534 7709 2534
rect 7961 1534 8011 2534
rect 9611 1534 9661 2534
rect 9913 1534 9963 2534
rect 11563 1534 11613 2534
rect 11865 1534 11915 2534
rect 13515 1534 13565 2534
rect 2905 290 2955 1290
rect 3755 290 3805 1290
rect 4057 290 4107 1290
rect 5707 290 5757 1290
rect 6009 290 6059 1290
rect 7659 290 7709 1290
rect 7961 290 8011 1290
rect 9611 290 9661 1290
rect 9913 290 9963 1290
rect 11563 290 11613 1290
rect 11865 290 11915 1290
rect 13515 290 13565 1290
<< metal2 >>
rect 99 -407 4879 -259
rect 5179 -407 5579 -210
rect 10078 -407 14858 -259
<< metal3 >>
rect 99 -407 4879 -16
rect 5179 -407 7379 -259
rect 7578 -407 9778 -89
rect 10078 -407 14858 -16
<< metal4 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 0 13600 254 18593
rect 14746 13600 15000 18593
rect 0 12410 254 13300
rect 14746 12410 15000 13300
rect 0 11240 254 12130
rect 14746 11240 15000 12130
rect 0 10874 254 10940
rect 14746 10874 15000 10940
rect 0 10218 100 10814
rect 14746 10218 14846 10814
rect 0 9922 254 10158
rect 14746 9922 15000 10158
rect 0 9266 116 9862
rect 14746 9266 14862 9862
rect 0 9140 254 9206
rect 14746 9140 15000 9206
rect 0 7910 254 8840
rect 14746 7910 15000 8840
rect 0 6940 254 7630
rect 14746 6940 15000 7630
rect 0 5970 254 6660
rect 14746 5970 15000 6660
rect 0 4760 254 5690
rect 14746 4760 15000 5690
rect 0 3550 254 4480
rect 14746 3550 15000 4480
rect 0 2580 254 3270
rect 14746 2580 15000 3270
rect 0 1370 254 2300
rect 14746 1370 15000 2300
rect 0 0 254 1090
rect 14746 0 15000 1090
<< metal5 >>
rect 0 34750 254 39593
rect 14746 34750 15000 39593
rect 7329 27458 7594 28780
rect 0 13600 254 18590
rect 14746 13600 15000 18590
rect 0 12430 254 13280
rect 14746 12430 15000 13280
rect 0 11260 254 12110
rect 14746 11260 15000 12110
rect 0 9140 254 10940
rect 14746 9140 15000 10940
rect 0 7930 254 8820
rect 14746 7930 15000 8820
rect 0 6960 254 7610
rect 14746 6960 15000 7610
rect 0 5990 254 6640
rect 14746 5990 15000 6640
rect 0 4780 254 5670
rect 14746 4780 15000 5670
rect 0 3570 254 4460
rect 14746 3570 15000 4460
rect 0 2600 254 3250
rect 14746 2600 15000 3250
rect 0 1390 254 2280
rect 14746 1390 15000 2280
rect 0 20 254 1070
rect 14746 20 15000 1070
use sky130_fd_io__top_power_hvc_wpadv2  sky130_fd_io__top_power_hvc_wpadv2_2 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602555073
transform 1 0 0 0 1 -407
box 0 0 15000 40000
use sky130_fd_io__overlay_vddio_hvc  sky130_fd_io__overlay_vddio_hvc_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1602555073
transform 1 0 0 0 1 -407
box 0 407 15000 40000
<< labels >>
flabel metal5 s 7329 27458 7594 28780 0 FreeSans 2000 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 127 37914 127 37914 3 FreeSans 520 0 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal4 s 14873 37914 14873 37914 3 FreeSans 520 180 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal2 s 10078 -407 14858 -259 2 FreeSans 2000 90 0 0 DRN_HVC
port 2 nsew power bidirectional
flabel metal2 s 99 -407 4879 -259 2 FreeSans 2000 90 0 0 SRC_BDY_HVC
port 4 nsew ground bidirectional
flabel metal3 s 7578 -407 9778 -89 0 FreeSans 2000 0 0 0 DRN_HVC
port 2 nsew power bidirectional
flabel metal3 s 10078 -407 14858 -16 0 FreeSans 2000 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal3 s 99 -407 4879 -16 0 FreeSans 2000 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal3 s 5179 -407 7379 -259 2 FreeSans 2000 90 0 0 SRC_BDY_HVC
port 4 nsew ground bidirectional
flabel metal5 s 14746 9140 15000 10940 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 14807 2600 15000 3250 3 FreeSans 520 180 0 0 VDDA
port 6 nsew power bidirectional
flabel metal5 s 14746 7930 15000 8820 3 FreeSans 520 180 0 0 VSSD
port 13 nsew ground bidirectional
flabel metal5 s 14746 11260 15000 12110 3 FreeSans 520 180 0 0 VSSIO_Q
port 14 nsew ground bidirectional
flabel metal5 s 14746 4780 15000 5670 3 FreeSans 520 180 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal5 s 14746 5990 15000 6640 3 FreeSans 520 180 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal5 s 14746 6961 15000 7610 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 14746 1390 15000 2280 3 FreeSans 520 180 0 0 VCCD
port 11 nsew power bidirectional
flabel metal5 s 14746 12430 15000 13280 3 FreeSans 520 180 0 0 VDDIO_Q
port 8 nsew power bidirectional
flabel metal5 s 14746 13600 15000 18590 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 14746 20 15000 1070 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal5 s 14746 3570 15000 4460 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 0 13600 254 18590 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 0 7930 254 8820 3 FreeSans 520 0 0 0 VSSD
port 13 nsew ground bidirectional
flabel metal5 s 0 11260 254 12110 3 FreeSans 520 0 0 0 VSSIO_Q
port 14 nsew ground bidirectional
flabel metal5 s 0 5990 254 6640 3 FreeSans 520 0 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal5 s 0 4780 254 5670 3 FreeSans 520 0 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal5 s 0 2600 193 3250 3 FreeSans 520 0 0 0 VDDA
port 6 nsew power bidirectional
flabel metal5 s 0 3570 254 4460 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal5 s 0 1390 254 2280 3 FreeSans 520 0 0 0 VCCD
port 11 nsew power bidirectional
flabel metal5 s 0 12430 254 13280 3 FreeSans 520 0 0 0 VDDIO_Q
port 8 nsew power bidirectional
flabel metal5 s 0 9140 254 10940 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 0 6961 254 7610 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal5 s 0 20 254 1070 3 FreeSans 520 0 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal4 s 14746 7910 15000 8840 3 FreeSans 520 180 0 0 VSSD
port 13 nsew ground bidirectional
flabel metal4 s 14807 2580 15000 3270 3 FreeSans 520 180 0 0 VDDA
port 6 nsew power bidirectional
flabel metal4 s 14746 11240 15000 12130 3 FreeSans 520 180 0 0 VSSIO_Q
port 14 nsew ground bidirectional
flabel metal4 s 14746 4760 15000 5690 3 FreeSans 520 180 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal4 s 14746 5970 15000 6660 3 FreeSans 520 180 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal4 s 14746 9922 15000 10158 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 14746 10874 15000 10940 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 14746 0 15000 1090 3 FreeSans 520 180 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal4 s 14746 3550 15000 4480 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 14746 9140 15000 9206 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 14746 6940 15000 7630 3 FreeSans 520 180 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 14746 12410 15000 13300 3 FreeSans 520 180 0 0 VDDIO_Q
port 8 nsew power bidirectional
flabel metal4 s 14746 1370 15000 2300 3 FreeSans 520 180 0 0 VCCD
port 11 nsew power bidirectional
flabel metal4 s 14746 9266 15000 9862 3 FreeSans 520 180 0 0 AMUXBUS_B
port 1 nsew signal bidirectional
flabel metal4 s 14746 34750 15000 39593 3 FreeSans 520 180 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal4 s 14746 10218 15000 10814 3 FreeSans 520 180 0 0 AMUXBUS_A
port 0 nsew signal bidirectional
flabel metal4 s 14746 13600 15000 18593 3 FreeSans 520 180 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 0 34750 254 39593 3 FreeSans 520 0 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal4 s 0 3550 254 4480 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 0 12410 254 13300 3 FreeSans 520 0 0 0 VDDIO_Q
port 8 nsew power bidirectional
flabel metal4 s 0 13600 254 18593 3 FreeSans 520 0 0 0 VDDIO
port 10 nsew power bidirectional
flabel metal4 s 0 1370 254 2300 3 FreeSans 520 0 0 0 VCCD
port 11 nsew power bidirectional
flabel metal4 s 0 9140 254 9206 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 5970 254 6660 3 FreeSans 520 0 0 0 VSWITCH
port 7 nsew power bidirectional
flabel metal4 s 0 0 254 1090 3 FreeSans 520 0 0 0 VCCHIB
port 9 nsew power bidirectional
flabel metal4 s 0 9922 254 10158 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 11240 254 12130 3 FreeSans 520 0 0 0 VSSIO_Q
port 14 nsew ground bidirectional
flabel metal4 s 0 4760 254 5690 3 FreeSans 520 0 0 0 VSSIO
port 12 nsew ground bidirectional
flabel metal4 s 0 2580 193 3270 3 FreeSans 520 0 0 0 VDDA
port 6 nsew power bidirectional
flabel metal4 s 0 10218 254 10814 3 FreeSans 520 0 0 0 AMUXBUS_A
port 0 nsew signal bidirectional
flabel metal4 s 0 10874 254 10940 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 6940 254 7630 3 FreeSans 520 0 0 0 VSSA
port 5 nsew ground bidirectional
flabel metal4 s 0 7910 254 8840 3 FreeSans 520 0 0 0 VSSD
port 13 nsew ground bidirectional
flabel metal4 s 0 9266 254 9862 3 FreeSans 520 0 0 0 AMUXBUS_B
port 1 nsew signal bidirectional
<< properties >>
string LEFclass PAD POWER
string FIXED_BBOX 0 0 15000 39593
<< end >>
