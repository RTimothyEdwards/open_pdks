magic
tech s8seal_ring
magscale 1 10
timestamp 1584558468
<< type81_51 >>
tri -14938 151666 0 152400 se
tri 0 151666 14938 152400 sw
tri -29732 149472 -14938 151666 se
rect -14938 149472 14938 151666
tri 14938 149472 29732 151666 sw
tri -44239 145838 -29732 149472 se
rect -29732 145838 29732 149472
tri 29732 145838 44239 149472 sw
tri -58321 140799 -44239 145838 se
rect -44239 140799 44239 145838
tri 44239 140799 58321 145838 sw
tri -71841 134405 -58321 140799 se
rect -58321 134405 58321 140799
tri 58321 134405 71841 140799 sw
tri -84669 126716 -71841 134405 se
rect -71841 126716 71841 134405
tri 71841 126716 84669 134405 sw
tri -96682 117807 -84669 126716 se
rect -84669 117807 84669 126716
tri 84669 117807 96682 126716 sw
tri -107763 107763 -96682 117807 se
rect -96682 107763 96682 117807
tri 96682 107763 107763 117807 sw
tri -117807 96682 -107763 107763 se
rect -107763 96682 107763 107763
tri 107763 96682 117807 107763 sw
tri -126716 84669 -117807 96682 se
rect -117807 84669 117807 96682
tri 117807 84669 126716 96682 sw
tri -134405 71841 -126716 84669 se
rect -126716 71841 126716 84669
tri 126716 71841 134405 84669 sw
tri -140799 58321 -134405 71841 se
rect -134405 58321 134405 71841
tri 134405 58321 140799 71841 sw
tri -145838 44239 -140799 58321 se
rect -140799 44239 140799 58321
tri 140799 44239 145838 58321 sw
tri -149472 29732 -145838 44239 se
rect -145838 29732 145838 44239
tri 145838 29732 149472 44239 sw
tri -151666 14938 -149472 29732 se
rect -149472 14938 149472 29732
tri 149472 14938 151666 29732 sw
tri -152400 0 -151666 14938 se
tri -152400 -14938 -151666 0 ne
rect -151666 -14938 151666 14938
tri 151666 0 152400 14938 sw
tri 151666 -14938 152400 0 nw
tri -151666 -29732 -149472 -14938 ne
rect -149472 -29732 149472 -14938
tri 149472 -29732 151666 -14938 nw
tri -149472 -44239 -145838 -29732 ne
rect -145838 -44239 145838 -29732
tri 145838 -44239 149472 -29732 nw
tri -145838 -58321 -140799 -44239 ne
rect -140799 -58321 140799 -44239
tri 140799 -58321 145838 -44239 nw
tri -140799 -71841 -134405 -58321 ne
rect -134405 -71841 134405 -58321
tri 134405 -71841 140799 -58321 nw
tri -134405 -84669 -126716 -71841 ne
rect -126716 -84669 126716 -71841
tri 126716 -84669 134405 -71841 nw
tri -126716 -96682 -117807 -84669 ne
rect -117807 -96682 117807 -84669
tri 117807 -96682 126716 -84669 nw
tri -117807 -107763 -107763 -96682 ne
rect -107763 -107763 107763 -96682
tri 107763 -107763 117807 -96682 nw
tri -107763 -117807 -96682 -107763 ne
rect -96682 -117807 96682 -107763
tri 96682 -117807 107763 -107763 nw
tri -96682 -126716 -84669 -117807 ne
rect -84669 -126716 84669 -117807
tri 84669 -126716 96682 -117807 nw
tri -84669 -134405 -71841 -126716 ne
rect -71841 -134405 71841 -126716
tri 71841 -134405 84669 -126716 nw
tri -71841 -140799 -58321 -134405 ne
rect -58321 -140799 58321 -134405
tri 58321 -140799 71841 -134405 nw
tri -58321 -145838 -44239 -140799 ne
rect -44239 -145838 44239 -140799
tri 44239 -145838 58321 -140799 nw
tri -44239 -149472 -29732 -145838 ne
rect -29732 -149472 29732 -145838
tri 29732 -149472 44239 -145838 nw
tri -29732 -151666 -14938 -149472 ne
rect -14938 -151666 14938 -149472
tri 14938 -151666 29732 -149472 nw
tri -14938 -152400 0 -151666 ne
tri 0 -152400 14938 -151666 nw
<< end >>
