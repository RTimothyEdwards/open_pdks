*
* spice test file for generating .prm files.
*
.lib /home/tim/projects/efabless/tech/XFAB/EFXH018D/libs.tech/models/lpmos/param.lib 3s
.lib /home/tim/projects/efabless/tech/XFAB/EFXH018D/libs.tech/models/lpmos/xh018.lib tm
*
.option TEMP=-5
*
* out1 - Output of Inverter to measure step response.
*
X0 out1 in1 GND GND ne L=0.18u W=0.8u
X1 out1 in1 VDD VDD pe L=0.18u W=1.0u
*
* out2 - Output of Inverter driven by out1 to determine slow-input effect.
*
X6 out2 out1 GND GND ne L=0.18u W=0.8u
X7 out2 out1 VDD VDD pe L=0.18u W=1.0u
*
* out3 - Output of a ne pulling up to determine dynamic-high resistance.
*
X2 out3 in2 VDD GND ne L=0.18u W=0.8u
*
* out4 - Output of a pe pulling down to determine dynamic-low resistance.
*
X3 out4 in3 GND VDD pe L=0.18u W=1.0u
*
* loading capacitors
*
C0 out1 GND 50f
C1 out2 GND 50f
C2 out3 GND 50f
C3 out4 GND 50f

VDD VDD 0 DC 1.98
* VGnd GND 0 DC 0
RGnd GND 0 0.01
Vmid mid 0 DC 0.9

Vin1 in1 0 0 pwl (0ns 0 0.1ns 1.98 40ns 1.98 40.1ns 0)
Vin2 in2 0 0 pwl (0ns 0 0.1ns 1.98)
Vin3 in3 0 5 pwl (0ns 1.98 0.1ns 0)

.ic V(out4)=1.98

.tran 0.01ns 80ns

.save all

.end
