magic
tech sky130A
magscale 1 2
timestamp 1602968705
<< error_p >>
rect 5750 2820 5758 2832
rect 5762 2786 5770 2820
rect 1886 2546 1916 2550
rect 1700 2540 1730 2544
rect 1730 2510 1734 2540
rect 1916 2516 1920 2546
rect 1692 2356 1722 2360
rect 1722 2326 1726 2356
rect 1896 2352 1926 2356
rect 1926 2322 1930 2352
rect 1694 2204 1724 2208
rect 1724 2174 1728 2204
rect 2216 2194 2286 2626
rect 3708 2524 3712 2558
rect 3928 2530 3942 2564
rect 4992 2490 5026 2492
rect 4992 2458 5026 2462
rect 5232 2458 5266 2462
rect 4374 2432 4408 2434
rect 5232 2428 5266 2432
rect 4522 2426 4556 2428
rect 5752 2418 5760 2430
rect 4374 2400 4408 2404
rect 4522 2394 4556 2396
rect 5764 2384 5772 2418
rect 2784 2238 2854 2374
rect 3700 2340 3704 2374
rect 3938 2336 3952 2370
rect 4538 2232 4572 2234
rect 3702 2188 3706 2222
rect 4538 2200 4572 2204
rect 5731 1620 5742 1631
rect 5768 1620 5779 1631
rect 5759 1557 5779 1607
rect 5809 1520 5829 1557
rect 5839 1520 5845 1557
rect 6229 1519 6232 1567
rect 6586 1503 6589 1551
rect 3240 1478 3256 1502
rect 6942 1500 6944 1547
rect 2406 1450 2440 1468
rect 3208 1454 3232 1470
rect 5720 1465 5731 1476
rect 5779 1465 5790 1476
rect 7415 1465 7417 1512
rect 2382 1410 2394 1444
rect 2406 1442 2440 1444
rect 2438 1414 2440 1442
rect 2406 1410 2440 1414
rect 2446 1410 2464 1444
rect 4867 1440 4945 1449
rect 5105 1436 5183 1444
rect 1936 1386 1948 1392
rect 1958 1386 1970 1392
rect 2406 1386 2440 1406
rect 1924 1368 1928 1380
rect 1936 1378 1970 1380
rect 1978 1368 1982 1380
rect 1924 1346 1928 1358
rect 1936 1346 1970 1348
rect 1978 1346 1982 1358
rect 1936 1334 1948 1340
rect 1958 1334 1970 1340
rect 4476 1324 4492 1330
rect 4494 1324 4510 1330
rect 3250 1284 3266 1308
rect 4460 1298 4466 1314
rect 4520 1298 4526 1314
rect 3902 1286 3936 1290
rect 4460 1280 4466 1296
rect 4520 1280 4526 1296
rect 3218 1260 3242 1276
rect 4476 1264 4492 1270
rect 4494 1264 4510 1270
rect 2420 1238 2454 1258
rect 2396 1200 2406 1234
rect 2420 1230 2454 1234
rect 2420 1200 2454 1204
rect 2464 1200 2478 1234
rect 1952 1192 1964 1198
rect 1940 1174 1942 1186
rect 1952 1184 1986 1186
rect 2420 1176 2454 1196
rect 1940 1152 1942 1164
rect 1952 1152 1986 1156
rect 1952 1140 1964 1148
rect 2498 666 2626 682
<< nwell >>
rect 5462 2652 6054 2988
rect 1620 2450 1984 2632
rect 3584 2466 4034 2634
rect 4300 2336 4618 2518
rect 4924 2394 5092 2576
rect 1714 1288 2032 1470
rect 2338 1346 2506 1528
rect 3132 1414 3302 1596
rect 5025 1330 5287 1700
rect 5588 1357 5929 1693
rect 7311 1307 7731 1732
<< nmos >>
rect 6229 1463 6285 1621
rect 7950 1405 7992 2994
<< scnmos >>
rect 6942 1444 6998 1602
<< scpmos >>
rect 7415 1409 7471 1567
<< varactor >>
rect 5731 1465 5779 1620
<< nmoslvt >>
rect 6586 1447 6642 1605
<< ndiff >>
rect 1674 2356 1744 2378
rect 1674 2326 1692 2356
rect 1722 2326 1744 2356
rect 1674 2306 1744 2326
rect 3620 2374 3754 2394
rect 3620 2340 3636 2374
rect 3670 2340 3700 2374
rect 3734 2340 3754 2374
rect 3620 2322 3754 2340
rect 5584 2322 5760 2496
rect 4514 2234 4604 2240
rect 4514 2200 4538 2234
rect 4572 2200 4604 2234
rect 4514 2196 4604 2200
rect 6176 1556 6229 1621
rect 6176 1519 6185 1556
rect 6221 1519 6229 1556
rect 6176 1463 6229 1519
rect 6285 1463 6348 1621
rect 6533 1540 6586 1605
rect 6533 1503 6542 1540
rect 6578 1503 6586 1540
rect 6533 1447 6586 1503
rect 6642 1447 6705 1605
rect 6889 1537 6942 1602
rect 6889 1500 6898 1537
rect 6934 1500 6942 1537
rect 6889 1444 6942 1500
rect 6998 1444 7061 1602
rect 7883 1405 7950 2994
rect 7992 1405 8098 2994
rect 1942 1186 2000 1192
rect 1942 1152 1952 1186
rect 1986 1152 2000 1186
rect 1942 1148 2000 1152
<< pdiff >>
rect 5582 2722 5758 2896
rect 1682 2540 1752 2562
rect 1682 2510 1700 2540
rect 1730 2510 1752 2540
rect 1682 2490 1752 2510
rect 3628 2558 3762 2578
rect 3628 2524 3644 2558
rect 3678 2524 3708 2558
rect 3742 2524 3762 2558
rect 3628 2506 3762 2524
rect 4498 2428 4582 2434
rect 4498 2394 4522 2428
rect 4556 2394 4582 2428
rect 4498 2388 4582 2394
rect 5105 1436 5183 1522
rect 1928 1380 1978 1386
rect 1928 1346 1936 1380
rect 1970 1346 1978 1380
rect 7362 1502 7415 1567
rect 7362 1465 7371 1502
rect 7407 1465 7415 1502
rect 7362 1409 7415 1465
rect 7471 1409 7534 1567
rect 1928 1340 1978 1346
<< ndiffc >>
rect 1692 2326 1722 2356
rect 3636 2340 3670 2374
rect 3700 2340 3734 2374
rect 4538 2200 4572 2234
rect 6185 1519 6221 1556
rect 6542 1503 6578 1540
rect 6898 1500 6934 1537
rect 1952 1152 1986 1186
<< pdiffc >>
rect 1700 2510 1730 2540
rect 3644 2524 3678 2558
rect 3708 2524 3742 2558
rect 4522 2394 4556 2428
rect 1936 1346 1970 1380
rect 7371 1465 7407 1502
<< psubdiff >>
rect 1872 2352 1950 2378
rect 1872 2322 1896 2352
rect 1926 2322 1950 2352
rect 1872 2298 1950 2322
rect 5204 2462 5294 2466
rect 3860 2370 3998 2398
rect 5204 2428 5232 2462
rect 5266 2428 5294 2462
rect 5204 2424 5294 2428
rect 3860 2336 3884 2370
rect 3918 2336 3938 2370
rect 3972 2336 3998 2370
rect 3860 2312 3998 2336
rect 5760 2418 5936 2496
rect 5760 2384 5764 2418
rect 5798 2384 5936 2418
rect 5760 2322 5936 2384
rect 4867 1440 4945 1526
rect 3184 1318 3250 1344
rect 3184 1284 3208 1318
rect 3242 1284 3250 1318
rect 3184 1276 3250 1284
rect 2406 1234 2464 1238
rect 2406 1200 2420 1234
rect 2454 1200 2464 1234
rect 2406 1196 2464 1200
rect 2458 666 2668 786
<< nsubdiff >>
rect 5758 2820 5934 2896
rect 5758 2786 5762 2820
rect 5796 2786 5934 2820
rect 5758 2722 5934 2786
rect 1862 2546 1940 2572
rect 1862 2516 1886 2546
rect 1916 2516 1940 2546
rect 1862 2492 1940 2516
rect 3848 2564 3986 2592
rect 3848 2530 3874 2564
rect 3908 2530 3928 2564
rect 3962 2530 3986 2564
rect 3848 2506 3986 2530
rect 4962 2492 5054 2498
rect 4962 2458 4992 2492
rect 5026 2458 5054 2492
rect 4962 2454 5054 2458
rect 4344 2434 4436 2440
rect 4344 2400 4374 2434
rect 4408 2400 4436 2434
rect 4344 2396 4436 2400
rect 5101 1637 5188 1662
rect 5101 1601 5129 1637
rect 5164 1601 5188 1637
rect 5101 1577 5188 1601
rect 3174 1512 3240 1538
rect 3174 1478 3198 1512
rect 3232 1478 3240 1512
rect 3174 1470 3240 1478
rect 2394 1444 2446 1450
rect 2394 1410 2406 1444
rect 2440 1410 2446 1444
rect 5681 1465 5731 1620
rect 5779 1557 5847 1620
rect 5779 1520 5809 1557
rect 5845 1520 5847 1557
rect 5779 1465 5847 1520
rect 2394 1406 2446 1410
rect 1764 1386 1846 1398
rect 1764 1352 1788 1386
rect 1822 1352 1846 1386
rect 1764 1340 1846 1352
rect 7621 1519 7691 1549
rect 7621 1482 7637 1519
rect 7673 1482 7691 1519
rect 7621 1457 7691 1482
<< psubdiffcont >>
rect 1896 2322 1926 2352
rect 5232 2428 5266 2462
rect 3884 2336 3918 2370
rect 3938 2336 3972 2370
rect 5764 2384 5798 2418
rect 3208 1284 3242 1318
rect 2420 1200 2454 1234
<< nsubdiffcont >>
rect 5762 2786 5796 2820
rect 1886 2516 1916 2546
rect 3874 2530 3908 2564
rect 3928 2530 3962 2564
rect 4992 2458 5026 2492
rect 4374 2400 4408 2434
rect 5129 1601 5164 1637
rect 3198 1478 3232 1512
rect 2406 1410 2440 1444
rect 5809 1520 5845 1557
rect 1788 1352 1822 1386
rect 7637 1482 7673 1519
<< poly >>
rect 7950 2994 7992 3045
rect 1676 2204 1746 2226
rect 1676 2174 1694 2204
rect 1724 2174 1746 2204
rect 3622 2222 3756 2242
rect 1676 2154 1746 2174
rect 3622 2188 3638 2222
rect 3672 2188 3702 2222
rect 3736 2188 3756 2222
rect 3622 2170 3756 2188
rect 5731 1620 5779 1665
rect 6229 1621 6285 1692
rect 5731 1420 5779 1465
rect 6586 1605 6642 1676
rect 6229 1417 6285 1463
rect 6942 1602 6998 1673
rect 4871 1402 4941 1412
rect 4871 1368 4887 1402
rect 4921 1368 4941 1402
rect 4871 1358 4941 1368
rect 5109 1397 5179 1407
rect 6586 1401 6642 1447
rect 7415 1567 7471 1638
rect 6942 1398 6998 1444
rect 5109 1363 5125 1397
rect 5159 1363 5179 1397
rect 7415 1363 7471 1409
rect 5109 1353 5179 1363
rect 7950 1351 7992 1405
rect 3886 1320 3956 1340
rect 3886 1286 3902 1320
rect 3936 1286 3956 1320
rect 3886 1280 3956 1286
rect 4466 1314 4520 1324
rect 4466 1280 4476 1314
rect 4510 1280 4520 1314
rect 4466 1270 4520 1280
rect 2529 635 2599 646
rect 2529 601 2545 635
rect 2579 601 2599 635
rect 2529 591 2599 601
<< polycont >>
rect 1694 2174 1724 2204
rect 3638 2188 3672 2222
rect 3702 2188 3736 2222
rect 4887 1368 4921 1402
rect 5125 1363 5159 1397
rect 3902 1286 3936 1320
rect 4476 1280 4510 1314
rect 2545 601 2579 635
<< xpolycontact >>
rect 2216 2194 2278 2626
rect 2784 2238 2854 2374
<< locali >>
rect 5762 2820 5796 2860
rect 5762 2752 5796 2786
rect 1848 2546 1952 2548
rect 1666 2540 1770 2542
rect 1666 2510 1700 2540
rect 1730 2510 1770 2540
rect 1848 2516 1886 2546
rect 1916 2516 1952 2546
rect 1848 2514 1952 2516
rect 1666 2508 1770 2510
rect 1658 2356 1762 2358
rect 1658 2326 1692 2356
rect 1722 2326 1762 2356
rect 1658 2324 1762 2326
rect 1860 2352 1964 2354
rect 1860 2322 1896 2352
rect 1926 2322 1964 2352
rect 1860 2320 1964 2322
rect 1660 2204 1764 2206
rect 1660 2174 1694 2204
rect 1724 2174 1764 2204
rect 3612 2524 3644 2558
rect 3678 2524 3708 2558
rect 3742 2524 3780 2558
rect 3838 2530 3874 2564
rect 3908 2530 3928 2564
rect 3962 2530 3996 2564
rect 4956 2458 4992 2492
rect 5026 2458 5060 2492
rect 4338 2400 4374 2434
rect 4408 2400 4442 2434
rect 5198 2428 5232 2462
rect 5266 2428 5302 2462
rect 4490 2394 4522 2428
rect 4556 2394 4594 2428
rect 5764 2418 5798 2454
rect 3604 2340 3636 2374
rect 3670 2340 3700 2374
rect 3734 2340 3772 2374
rect 3850 2336 3884 2370
rect 3918 2336 3938 2370
rect 3972 2336 4008 2370
rect 5764 2348 5798 2384
rect 3606 2188 3638 2222
rect 3672 2188 3702 2222
rect 3736 2188 3774 2222
rect 4506 2200 4538 2234
rect 4572 2200 4610 2234
rect 1660 2172 1764 2174
rect 5088 1637 5220 1638
rect 5088 1601 5129 1637
rect 5164 1601 5220 1637
rect 5809 1557 5845 1593
rect 3162 1478 3198 1512
rect 3232 1478 3266 1512
rect 5809 1487 5845 1520
rect 6185 1556 6221 1587
rect 6185 1487 6221 1519
rect 6542 1540 6578 1571
rect 6542 1471 6578 1503
rect 6898 1537 6934 1568
rect 6898 1468 6934 1500
rect 7371 1502 7407 1533
rect 2370 1410 2406 1444
rect 2440 1410 2474 1444
rect 7371 1433 7407 1465
rect 7637 1519 7673 1553
rect 7637 1441 7673 1482
rect 1752 1352 1788 1386
rect 1822 1352 1856 1386
rect 1904 1346 1936 1380
rect 1970 1346 2008 1380
rect 4855 1368 4887 1402
rect 4921 1368 4959 1402
rect 5093 1363 5125 1397
rect 5159 1363 5197 1397
rect 3174 1284 3208 1318
rect 3242 1284 3278 1318
rect 3870 1286 3902 1320
rect 3936 1286 3974 1320
rect 4444 1280 4476 1314
rect 4510 1280 4548 1314
rect 2386 1200 2420 1234
rect 2454 1200 2490 1234
rect 1920 1152 1952 1186
rect 1986 1152 2024 1186
rect 2513 601 2545 635
rect 2579 601 2617 635
<< labels >>
flabel comment s 408 552 408 552 0 FreeSans 560 0 0 0 Not implemented
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Licon
flabel comment s 1740 2062 1740 2068 0 FreeSans 560 0 0 0 licon.1
flabel comment s 2326 2076 2326 2082 0 FreeSans 560 0 0 0 licon.1b
flabel comment s 2894 2094 2894 2100 0 FreeSans 560 0 0 0 licon.1c
flabel comment s 3834 2046 3834 2052 0 FreeSans 560 0 0 0 licon.2
flabel comment s 476 334 476 334 0 FreeSans 560 0 0 0 licon 2b, 2c, 2d
flabel comment s 4902 2084 4902 2090 0 FreeSans 560 0 0 0 licon.5a
flabel comment s 5816 2128 5816 2134 0 FreeSans 560 0 0 0 licon.5b
flabel comment s 2316 1036 2316 1042 0 FreeSans 560 0 0 0 licon.5c
flabel comment s 3250 1108 3250 1108 0 FreeSans 560 0 0 0 licon.7
flabel comment s 3926 1108 3926 1108 0 FreeSans 560 0 0 0 licon.8
flabel comment s 4460 1094 4460 1094 0 FreeSans 560 0 0 0 licon.8a
flabel comment s 5067 1151 5067 1151 0 FreeSans 560 0 0 0 licon.9
flabel comment s 5767 1227 5767 1227 0 FreeSans 560 0 0 0 licon.10
flabel comment s 6300 1265 6300 1265 0 FreeSans 560 0 0 0 licon.11
flabel comment s 482 145 482 145 0 FreeSans 560 0 0 0 licon 11c, 11d
flabel comment s 6989 1257 6989 1257 0 FreeSans 560 0 0 0 licon.11a
flabel comment s 7977 1246 7977 1246 0 FreeSans 560 0 0 0 licon.12
flabel comment s 8055 3214 8055 3214 0 FreeSans 560 0 0 0 Not implemented
flabel comment s 7526 1216 7526 1216 0 FreeSans 560 0 0 0 licon.11b
flabel comment s 2632 390 2632 390 0 FreeSans 560 0 0 0 licon.14
flabel comment s 2628 515 2628 515 0 FreeSans 560 0 0 0 licon.13
flabel comment s 478 -4 478 -4 0 FreeSans 560 0 0 0 licon.16
flabel comment s 473 1576 479 1576 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s 399 1412 399 1412 0 FreeSans 560 0 0 0 licon.3
flabel comment s 409 1292 409 1292 0 FreeSans 560 0 0 0 licon.4
flabel comment s 409 1170 409 1170 0 FreeSans 560 0 0 0 licon.6
flabel comment s 395 1020 395 1020 0 FreeSans 560 0 0 0 licon.15
flabel comment s 425 912 425 912 0 FreeSans 560 0 0 0 licon.17
flabel comment s 440 789 440 789 0 FreeSans 560 0 0 0 licon.18
flabel comment s 454 -272 454 -272 0 FreeSans 560 0 0 0 Do not understand
flabel comment s 514 -421 514 -421 0 FreeSans 560 0 0 0 licon.19
<< end >>
