MACRO sky130_fd_io__top_xres4v2
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_xres4v2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY R90 ;
  PIN PAD_A_ESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.245 0.000 18.910 0.565 ;
    END
    PORT
      LAYER met2 ;
        RECT 17.245 0.000 18.910 0.565 ;
    END
  END PAD_A_ESD_H
  PIN XRES_H_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.935 0.000 29.665 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.935 0.000 29.665 0.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170 10.610 28.900 13.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170 10.610 29.050 10.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170 10.910 28.900 14.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.170 10.145 28.635 10.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.335 10.445 29.215 10.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.635 9.845 29.665 10.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.900 10.145 29.665 10.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.935 0.000 29.665 9.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.935 4.005 29.665 10.145 ;
    END
  END XRES_H_N
  PIN FILT_IN_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.075 0.000 21.225 1.410 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.075 0.000 21.225 1.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075 3.410 21.225 8.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075 6.820 21.375 6.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075 6.970 21.525 7.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075 7.120 21.675 7.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.075 7.150 21.060 8.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.225 7.150 21.705 7.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.375 7.300 21.855 7.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.525 7.450 22.005 7.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.675 7.600 22.155 7.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.825 7.750 22.305 7.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.060 8.135 22.970 8.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.225 6.670 22.690 8.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.340 8.415 24.050 9.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.575 8.500 23.055 8.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.725 8.650 23.205 8.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.875 8.800 23.355 8.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 8.950 23.505 9.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.175 9.100 23.655 9.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.325 9.250 23.805 9.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 9.495 24.050 9.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.690 8.135 22.970 8.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.720 9.645 24.050 9.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 9.495 24.050 9.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 9.980 24.050 12.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.970 8.415 24.050 9.495 ;
    END
  END FILT_IN_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.400 0.000 8.920 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 8.425 0.000 8.895 0.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775 17.410 7.295 31.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775 17.410 7.400 17.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775 17.515 7.295 17.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775 17.620 7.295 31.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775 31.400 7.400 31.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775 31.505 7.150 31.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.775 16.895 7.290 17.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.925 31.505 7.505 31.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.150 31.880 8.595 32.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.290 16.445 8.330 17.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.290 16.895 7.870 17.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.295 17.045 7.870 17.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.295 31.295 7.880 31.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.375 31.955 7.955 32.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 16.745 8.020 16.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.525 32.105 8.105 32.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.675 32.255 8.255 32.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.740 15.995 8.920 16.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.865 32.595 9.180 33.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.870 16.585 8.330 17.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.880 31.880 8.595 32.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.890 16.295 8.470 16.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.125 32.705 8.705 32.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.190 15.785 8.920 15.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.275 32.855 8.855 33.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.330 15.995 8.920 16.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.400 0.000 8.920 15.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.400 1.135 8.920 15.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.450 33.180 9.395 33.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.595 32.595 9.180 33.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.815 33.395 22.275 33.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.970 33.700 21.970 34.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.115 33.695 22.275 33.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.180 33.180 9.395 33.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.395 33.995 22.275 34.125 ;
    END
  END ENABLE_VDDIO
  PIN TIE_WEAK_HI_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.190 0.000 73.260 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 72.215 0.000 73.235 0.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860 71.930 65.990 93.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860 71.930 66.310 72.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860 72.080 66.160 72.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860 72.400 65.990 94.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.860 70.750 66.040 71.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.140 71.650 66.590 71.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.290 71.500 66.740 71.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.440 71.350 66.890 71.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.590 71.200 67.040 71.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.990 72.210 66.180 72.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.040 69.400 68.355 71.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.040 70.750 67.490 70.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.180 71.000 67.390 72.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.190 70.600 67.640 70.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.340 70.450 67.790 70.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.490 70.300 67.940 70.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 70.150 68.090 70.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.940 69.850 68.390 70.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.090 69.700 68.540 69.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390 68.535 69.305 69.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390 69.400 68.840 69.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.390 70.035 68.355 71.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.540 69.250 68.990 69.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.690 69.100 69.140 69.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.990 68.800 69.440 68.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.255 67.600 70.590 68.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 68.500 69.740 68.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.355 69.085 69.305 70.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.440 68.350 69.890 68.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.590 68.200 70.040 68.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 68.050 70.190 68.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190 66.200 72.190 67.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.190 67.600 70.640 67.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.305 67.800 70.590 69.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 67.450 70.790 67.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.490 67.300 70.940 67.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.640 67.150 71.090 67.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.790 67.000 71.240 67.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.940 66.850 71.390 67.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.090 66.700 71.540 66.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.240 66.550 71.690 66.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.390 66.400 71.840 66.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.590 64.600 73.925 66.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.590 66.200 72.190 67.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.840 65.950 72.290 66.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.990 65.800 72.440 65.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.140 65.650 72.590 65.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.290 65.500 72.740 65.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.440 65.350 72.890 65.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.590 65.200 73.040 65.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.740 65.050 73.190 65.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.890 64.900 73.340 65.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 0.000 73.260 49.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 0.725 73.260 49.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 49.470 73.925 64.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 49.620 73.560 49.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 49.770 73.710 49.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 49.985 73.925 64.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 64.465 73.925 64.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 64.465 73.925 66.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 64.530 73.795 64.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 64.595 73.790 64.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.260 49.320 73.925 49.985 ;
    END
  END TIE_WEAK_HI_H
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.285 0.000 12.545 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 12.285 0.000 12.545 0.330 ;
    END
  END ENABLE_H
  PIN PULLUP_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.555 0.000 15.135 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 14.555 0.000 15.135 0.330 ;
    END
  END PULLUP_H
  PIN EN_VDDIO_SIG_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.360 0.000 22.660 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.360 0.000 22.660 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 4.250 10.375 4.580 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.965 9.200 10.535 9.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.005 3.905 10.350 4.250 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.165 9.400 10.865 9.730 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.210 4.045 10.510 4.115 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.295 9.460 10.595 9.530 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.335 9.200 10.535 9.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.350 3.575 10.930 3.930 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.365 9.530 10.665 9.600 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.375 3.930 10.695 4.250 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.420 3.835 10.720 3.905 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.490 3.765 10.790 3.835 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.495 9.730 11.125 10.100 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.535 9.400 10.865 9.730 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.575 9.740 10.875 9.810 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.645 9.810 10.945 9.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 26.610 11.125 27.300 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 26.825 11.125 27.085 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 27.085 10.910 28.005 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 27.085 11.055 27.155 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 27.155 10.985 27.225 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 27.295 10.910 27.300 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 27.300 10.910 27.935 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 28.005 11.125 28.625 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 28.075 11.050 28.145 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 28.150 11.125 28.410 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.650 28.410 10.865 28.625 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.655 26.820 11.125 26.825 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.680 3.435 15.245 3.575 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.680 3.575 15.025 3.645 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.695 3.695 10.930 3.930 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.715 9.880 11.015 9.950 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.720 28.410 11.125 28.480 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.725 26.750 11.125 26.820 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.790 28.480 11.125 28.550 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.820 3.435 14.885 3.695 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 10.045 11.125 10.100 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 10.100 11.125 26.610 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 28.150 11.125 31.140 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 28.620 11.125 28.625 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 28.625 11.125 31.085 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 31.140 11.270 31.455 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 31.195 11.125 31.455 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 9.730 11.125 9.990 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.865 9.990 11.125 27.085 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.910 27.085 11.125 27.300 ;
    END
    PORT
      LAYER met2 ;
        RECT 10.910 27.935 11.125 28.150 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.005 31.265 11.305 31.335 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.125 31.085 11.270 31.230 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.125 31.455 11.520 31.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.260 31.480 11.520 36.020 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.260 31.535 11.520 31.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.260 36.020 12.150 36.280 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.270 31.230 11.495 31.455 ;
    END
    PORT
      LAYER met2 ;
        RECT 11.495 31.455 11.520 31.480 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.775 3.695 15.245 3.795 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.875 3.795 15.515 4.065 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.885 3.435 15.245 3.795 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.985 3.835 15.285 3.905 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.055 3.905 15.355 3.975 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.145 4.065 15.885 4.435 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.245 3.795 15.515 4.065 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.265 4.115 15.565 4.185 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.335 4.185 15.635 4.255 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.405 4.255 15.705 4.325 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.515 4.065 15.885 4.435 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.515 4.435 15.995 4.805 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.615 4.465 15.915 4.535 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.695 4.545 28.765 4.615 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.765 4.615 28.835 4.685 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.885 4.435 15.995 4.545 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.885 4.755 28.975 4.805 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.060 4.245 22.660 4.545 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.065 4.540 22.940 4.545 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.135 4.470 22.870 4.540 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.205 4.400 22.800 4.470 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.345 4.260 22.660 4.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.350 4.255 22.660 4.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.360 0.000 22.660 4.245 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.360 1.170 22.660 4.805 ;
    END
    PORT
      LAYER met2 ;
        RECT 22.660 4.260 22.945 4.545 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.655 4.805 29.120 4.900 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.750 4.900 29.450 5.230 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.765 4.545 29.120 4.900 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.865 4.945 29.165 5.015 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.935 5.015 29.235 5.085 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.005 5.085 29.305 5.155 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.080 5.230 29.580 5.470 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.120 4.900 29.450 5.230 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320 10.975 29.770 11.165 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320 11.085 29.400 11.165 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320 5.360 29.580 11.030 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320 5.415 29.580 5.470 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320 5.470 29.580 10.975 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.400 11.165 30.030 11.535 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.450 5.230 29.580 5.360 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.530 11.225 29.830 11.295 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.580 10.975 29.770 11.165 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.600 11.295 29.900 11.365 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770 11.165 30.030 11.425 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770 11.425 30.030 15.700 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770 11.480 30.030 11.535 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770 11.535 30.030 15.645 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770 15.700 30.365 15.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.770 15.755 29.995 15.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.840 15.755 30.140 15.825 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.910 15.825 30.210 15.895 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.995 15.980 30.625 16.350 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.030 15.645 30.365 15.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.120 16.035 30.420 16.105 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.190 16.105 30.490 16.175 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.365 15.980 30.625 16.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.365 16.240 30.625 16.350 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.365 16.350 30.625 20.495 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 4.250 10.005 4.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 4.520 10.050 4.575 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 4.520 9.995 8.915 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 4.575 9.995 4.630 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 4.630 9.995 8.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 8.915 10.335 9.200 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.735 8.970 9.965 9.200 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.790 4.465 10.105 4.520 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.805 8.970 10.105 9.040 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.860 4.395 10.160 4.465 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.875 9.040 10.175 9.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.930 4.325 10.230 4.395 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.965 9.200 10.165 9.400 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.995 8.860 10.335 9.200 ;
    END
  END EN_VDDIO_SIG_H
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.580 0.000 28.230 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.580 0.000 28.230 0.330 ;
    END
  END TIE_LO_ESD
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.505 0.000 31.155 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 30.505 0.000 31.155 0.330 ;
    END
  END TIE_HI_ESD
  PIN DISABLE_PULLUP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.760 0.000 33.020 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 32.760 0.000 33.020 0.330 ;
    END
  END DISABLE_PULLUP_H
  PIN INP_SEL_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.905 0.000 25.135 9.975 ;
    END
  END INP_SEL_H
  PIN VSSIO
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
  END VSSIO
  PIN VSSA
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 1.270 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 1.270 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
  END VSSD
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 1.270 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 1.270 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
  END VDDIO
  PIN VSWITCH
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
  END VSWITCH
  PIN VDDA
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
  END VCCHIB
  PIN VSSIO_Q
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
  END VSSIO_Q
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 17.250 108.455 54.435 164.285 ;
    END
  END PAD
  OBS
      LAYER nwell ;
        RECT -0.515 168.515 75.620 170.210 ;
        RECT -0.515 146.690 1.675 168.515 ;
        RECT 73.095 146.690 75.620 168.515 ;
        RECT -0.515 144.880 75.620 146.690 ;
      LAYER pwell ;
        RECT -0.290 140.685 75.290 144.565 ;
      LAYER nwell ;
        RECT -0.330 130.665 75.330 140.380 ;
      LAYER pwell ;
        RECT -0.130 129.315 41.750 130.355 ;
        RECT 61.910 129.315 75.130 130.355 ;
        RECT -0.130 124.135 75.130 129.315 ;
        RECT -0.130 102.525 1.435 124.135 ;
        RECT 73.560 102.525 75.130 124.135 ;
        RECT -0.130 99.230 75.130 102.525 ;
        RECT -0.130 97.995 58.470 99.230 ;
        RECT 71.930 97.995 75.130 99.230 ;
        RECT -0.130 96.735 75.130 97.995 ;
        RECT -0.130 96.730 58.470 96.735 ;
      LAYER li1 ;
        RECT 0.000 144.435 75.000 199.220 ;
        RECT -0.160 140.815 75.160 144.435 ;
        RECT 0.000 130.225 75.000 140.815 ;
        RECT -0.265 101.395 75.000 130.225 ;
        RECT 0.000 0.185 75.000 101.395 ;
      LAYER met1 ;
        RECT 0.000 170.090 75.000 199.210 ;
        RECT -0.145 131.275 75.145 170.090 ;
        RECT 0.000 130.220 75.000 131.275 ;
        RECT -0.145 95.895 75.145 130.220 ;
        RECT 0.000 10.255 75.000 95.895 ;
        RECT 0.000 0.610 24.625 10.255 ;
        RECT 0.000 0.185 12.005 0.610 ;
        RECT 12.825 0.185 14.275 0.610 ;
        RECT 15.415 0.185 22.080 0.610 ;
        RECT 22.940 0.185 24.625 0.610 ;
        RECT 25.415 0.610 75.000 10.255 ;
        RECT 25.415 0.185 27.300 0.610 ;
        RECT 28.510 0.185 30.225 0.610 ;
        RECT 31.435 0.185 32.480 0.610 ;
        RECT 33.300 0.185 75.000 0.610 ;
      LAYER met2 ;
        RECT 0.340 36.560 74.915 199.210 ;
        RECT 0.340 31.870 10.980 36.560 ;
        RECT 12.430 35.740 74.915 36.560 ;
        RECT 0.340 31.735 10.845 31.870 ;
        RECT 0.340 28.905 10.585 31.735 ;
        RECT 11.800 31.175 74.915 35.740 ;
        RECT 11.775 30.950 74.915 31.175 ;
        RECT 11.550 30.805 74.915 30.950 ;
        RECT 0.340 26.330 10.370 28.905 ;
        RECT 11.405 27.655 74.915 30.805 ;
        RECT 11.190 27.580 74.915 27.655 ;
        RECT 0.340 10.380 10.585 26.330 ;
        RECT 11.405 20.775 74.915 27.580 ;
        RECT 11.405 16.630 30.085 20.775 ;
        RECT 11.405 16.260 29.715 16.630 ;
        RECT 11.405 11.815 29.490 16.260 ;
        RECT 30.905 15.700 74.915 20.775 ;
        RECT 30.645 15.365 74.915 15.700 ;
        RECT 11.405 11.445 29.120 11.815 ;
        RECT 0.340 10.010 10.215 10.380 ;
        RECT 0.340 9.680 9.885 10.010 ;
        RECT 0.340 9.480 9.685 9.680 ;
        RECT 0.340 3.970 9.455 9.480 ;
        RECT 11.405 9.450 29.040 11.445 ;
        RECT 30.310 10.885 74.915 15.365 ;
        RECT 30.050 10.695 74.915 10.885 ;
        RECT 11.145 9.120 29.040 9.450 ;
        RECT 10.815 8.920 29.040 9.120 ;
        RECT 10.615 8.580 29.040 8.920 ;
        RECT 10.275 5.750 29.040 8.580 ;
        RECT 10.275 5.510 28.800 5.750 ;
        RECT 10.275 5.180 28.470 5.510 ;
        RECT 10.275 5.085 28.375 5.180 ;
        RECT 10.275 4.860 15.235 5.085 ;
        RECT 29.860 4.950 74.915 10.695 ;
        RECT 10.655 4.715 15.235 4.860 ;
        RECT 10.655 4.530 14.865 4.715 ;
        RECT 29.730 4.620 74.915 4.950 ;
        RECT 10.975 4.345 14.865 4.530 ;
        RECT 10.975 4.210 14.595 4.345 ;
        RECT 29.400 4.265 74.915 4.620 ;
        RECT 11.210 4.075 14.595 4.210 ;
        RECT 16.275 4.155 21.780 4.265 ;
        RECT 11.210 3.975 14.495 4.075 ;
        RECT 0.340 3.625 9.725 3.970 ;
        RECT 16.165 3.965 21.780 4.155 ;
        RECT 23.225 3.980 74.915 4.265 ;
        RECT 16.165 3.785 22.080 3.965 ;
        RECT 0.340 3.295 10.070 3.625 ;
        RECT 15.795 3.515 22.080 3.785 ;
        RECT 0.340 3.155 10.400 3.295 ;
        RECT 15.525 3.155 22.080 3.515 ;
        RECT 0.340 1.690 22.080 3.155 ;
        RECT 0.340 0.845 19.795 1.690 ;
        RECT 0.340 0.610 16.965 0.845 ;
        RECT 0.340 0.000 8.145 0.610 ;
        RECT 9.175 0.000 12.005 0.610 ;
        RECT 12.825 0.000 14.275 0.610 ;
        RECT 15.415 0.000 16.965 0.610 ;
        RECT 19.190 0.000 19.795 0.845 ;
        RECT 21.505 0.000 22.080 1.690 ;
        RECT 22.940 0.610 74.915 3.980 ;
        RECT 22.940 0.000 27.300 0.610 ;
        RECT 28.510 0.000 28.655 0.610 ;
        RECT 29.945 0.000 30.225 0.610 ;
        RECT 31.435 0.000 32.480 0.610 ;
        RECT 33.300 0.000 71.935 0.610 ;
        RECT 73.515 0.000 74.915 0.610 ;
      LAYER met3 ;
        RECT 0.965 95.045 74.700 200.000 ;
        RECT 0.965 70.350 64.460 95.045 ;
        RECT 66.390 72.800 74.700 95.045 ;
        RECT 66.580 72.610 74.700 72.800 ;
        RECT 67.790 71.400 74.700 72.610 ;
        RECT 68.755 70.435 74.700 71.400 ;
        RECT 0.965 69.000 65.640 70.350 ;
        RECT 69.705 69.485 74.700 70.435 ;
        RECT 0.965 68.135 66.990 69.000 ;
        RECT 70.990 68.200 74.700 69.485 ;
        RECT 0.965 67.200 67.855 68.135 ;
        RECT 0.965 65.800 68.790 67.200 ;
        RECT 72.590 66.600 74.700 68.200 ;
        RECT 0.965 64.200 70.190 65.800 ;
        RECT 0.965 34.525 71.790 64.200 ;
        RECT 74.325 48.920 74.700 66.600 ;
        RECT 0.965 34.100 8.570 34.525 ;
        RECT 0.965 33.580 8.050 34.100 ;
        RECT 0.965 32.995 7.465 33.580 ;
        RECT 22.675 32.995 71.790 34.525 ;
        RECT 0.965 32.280 6.750 32.995 ;
        RECT 9.795 32.780 71.790 32.995 ;
        RECT 0.965 16.495 6.375 32.280 ;
        RECT 9.580 32.195 71.790 32.780 ;
        RECT 8.995 31.480 71.790 32.195 ;
        RECT 8.280 30.895 71.790 31.480 ;
        RECT 7.695 18.020 71.790 30.895 ;
        RECT 8.270 17.445 71.790 18.020 ;
        RECT 8.730 16.985 71.790 17.445 ;
        RECT 0.965 16.045 6.890 16.495 ;
        RECT 0.965 15.595 7.340 16.045 ;
        RECT 0.965 15.385 7.790 15.595 ;
        RECT 0.965 0.565 8.000 15.385 ;
        RECT 9.320 15.170 71.790 16.985 ;
        RECT 9.320 12.665 27.770 15.170 ;
        RECT 9.320 10.380 22.505 12.665 ;
        RECT 9.320 8.815 20.940 10.380 ;
        RECT 24.450 9.745 27.770 12.665 ;
        RECT 29.300 11.310 71.790 15.170 ;
        RECT 24.450 9.445 28.235 9.745 ;
        RECT 9.320 8.535 20.660 8.815 ;
        RECT 9.320 3.010 19.675 8.535 ;
        RECT 24.450 8.015 28.535 9.445 ;
        RECT 23.370 7.735 28.535 8.015 ;
        RECT 23.090 6.270 28.535 7.735 ;
        RECT 21.625 3.010 28.535 6.270 ;
        RECT 9.320 1.810 28.535 3.010 ;
        RECT 9.320 0.965 19.675 1.810 ;
        RECT 9.320 0.565 16.845 0.965 ;
        RECT 19.310 0.565 19.675 0.965 ;
        RECT 21.625 0.565 28.535 1.810 ;
        RECT 30.065 0.565 71.790 11.310 ;
        RECT 73.660 0.565 74.700 48.920 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 165.885 75.000 174.185 ;
        RECT 0.000 106.855 15.650 165.885 ;
        RECT 56.035 106.855 75.000 165.885 ;
        RECT 0.000 96.585 75.000 106.855 ;
        RECT 2.870 18.285 72.130 96.585 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__top_xres4v2
END LIBRARY

