* Power pads library (sky130 power pads + overlays)
* Includes corner and fill cell subcircuits

.SUBCKT sky130_ef_io__vdda_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vdda_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vddio_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vddio_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vccd_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vccd_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vssa_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vssa_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vssio_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vssio_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vssd_hvc_pad
+ amuxbus_a amuxbus_b drn_hvc src_bdy_hvc
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__vssd_lvc_pad
+ amuxbus_a amuxbus_b drn_lvc1 drn_lvc2 src_bdy_lvc1 src_bdy_lvc2
+ bdy2_b2b vssi
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__corner_pad
+ amuxbus_a amuxbus_b 
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__com_bus_slice
+ amuxbus_a amuxbus_b
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__com_bus_slice_1um
+ amuxbus_a amuxbus_b
+ vssa vdda vswitch vddio_q vcchib vddio vccd vssio vssd vssio_q
.ENDS

.SUBCKT sky130_ef_io__gpiov2_pad
+ in_h pad_a_noesd_h pad_a_esd_0_h pad_a_esd_1_h
+ pad dm<2> dm<1> dm<0> hld_h_n in inp_dis ib_mode_sel enable_h enable_vdda_h
+ enable_inp_h oe_n tie_hi_esd tie_lo_esd slow vtrip_sel hld_ovr
+ analog_en analog_sel enable_vddio enable_vswitch_h analog_pol out
+ amuxbus_a amuxbus_b vssa vdda vswitch vddio_q vcchib vddio vccd vssio
+ vssd vssio_q
.ENDS
