magic
tech s8seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
tri 410 2269 470 2294 se
tri 470 2269 495 2294 sw
tri 410 2184 495 2269 ne
tri 495 2184 580 2269 sw
tri 495 2099 580 2184 ne
tri 580 2099 665 2184 sw
tri 580 2014 665 2099 ne
tri 665 2014 750 2099 sw
tri 665 1929 750 2014 ne
tri 750 1929 835 2014 sw
tri 750 1844 835 1929 ne
tri 835 1844 920 1929 sw
tri 835 1759 920 1844 ne
tri 920 1759 1005 1844 sw
tri 920 1674 1005 1759 ne
tri 1005 1674 1090 1759 sw
tri 1005 1589 1090 1674 ne
tri 1090 1589 1175 1674 sw
tri 1090 1504 1175 1589 ne
tri 1175 1504 1260 1589 sw
tri 1175 1419 1260 1504 ne
tri 1260 1419 1345 1504 sw
tri 1260 1334 1345 1419 ne
tri 1345 1334 1430 1419 sw
tri 1345 1249 1430 1334 ne
tri 1430 1249 1515 1334 sw
tri 1430 1164 1515 1249 ne
tri 1515 1164 1600 1249 sw
tri 1515 1079 1600 1164 ne
tri 1600 1079 1685 1164 sw
tri 1600 994 1685 1079 ne
tri 1685 994 1770 1079 sw
tri 1685 909 1770 994 ne
tri 1770 909 1855 994 sw
tri 1770 824 1855 909 ne
tri 1855 824 1940 909 sw
tri 1855 739 1940 824 ne
tri 1940 739 2025 824 sw
tri 1940 654 2025 739 ne
tri 2025 654 2110 739 sw
tri 2025 569 2110 654 ne
tri 2110 569 2195 654 sw
tri 2110 484 2195 569 ne
tri 2195 484 2280 569 sw
tri 2195 410 2269 484 ne
rect 2269 470 2280 484
tri 2280 470 2294 484 sw
rect 2269 410 51200 470
<< end >>
