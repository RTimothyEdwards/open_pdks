magic
tech sky130seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
tri 650 2369 710 2394 se
tri 710 2369 735 2394 sw
tri 650 2284 735 2369 ne
tri 735 2284 820 2369 sw
tri 735 2199 820 2284 ne
tri 820 2199 905 2284 sw
tri 820 2114 905 2199 ne
tri 905 2114 990 2199 sw
tri 905 2029 990 2114 ne
tri 990 2029 1075 2114 sw
tri 990 1944 1075 2029 ne
tri 1075 1944 1160 2029 sw
tri 1075 1859 1160 1944 ne
tri 1160 1859 1245 1944 sw
tri 1160 1774 1245 1859 ne
tri 1245 1774 1330 1859 sw
tri 1245 1689 1330 1774 ne
tri 1330 1689 1415 1774 sw
tri 1330 1604 1415 1689 ne
tri 1415 1604 1500 1689 sw
tri 1415 1519 1500 1604 ne
tri 1500 1519 1585 1604 sw
tri 1500 1434 1585 1519 ne
tri 1585 1434 1670 1519 sw
tri 1585 1349 1670 1434 ne
tri 1670 1349 1755 1434 sw
tri 1670 1264 1755 1349 ne
tri 1755 1264 1840 1349 sw
tri 1755 1179 1840 1264 ne
tri 1840 1179 1925 1264 sw
tri 1840 1094 1925 1179 ne
tri 1925 1094 2010 1179 sw
tri 1925 1009 2010 1094 ne
tri 2010 1009 2095 1094 sw
tri 2010 924 2095 1009 ne
tri 2095 924 2180 1009 sw
tri 2095 839 2180 924 ne
tri 2180 839 2265 924 sw
tri 2180 754 2265 839 ne
tri 2265 754 2350 839 sw
tri 2265 669 2350 754 ne
tri 2350 710 2394 754 sw
rect 2350 669 51200 710
tri 2350 650 2369 669 ne
rect 2369 650 51200 669
<< end >>
