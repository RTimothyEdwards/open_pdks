VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;

SITE unithd
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE  0.460 BY 2.720 ;
END unithd

LAYER li1
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH 0.46 0.34 ;
    OFFSET 0.23 0.17 ;

    WIDTH    0.170 ;                    # LI 1
    # SPACING  0.170 ;                    # LI 2
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0 0.170000 ;
    AREA 0.0561 ;                       # LI 6
    THICKNESS 0.10 ; 

    RESISTANCE RPERSQ 12.2 ;

    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 75.0 ) ( 0.0125 75.0 ) ( 0.0225 85.125 ) ( 22.5 10200.0 ) ) ;


END li1

LAYER mcon
  TYPE CUT ;
  WIDTH   0.17 ;		# Mcon 1
  SPACING 0.19 ;		# Mcon 2
  ENCLOSURE BELOW 0.0 0.0 ;	# Mcon 4
  ENCLOSURE ABOVE 0.030 0.060 ; # Met1 4 / Met1 5

  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC
  ANTENNADIFFAREARATIO PWL ( ( 0.0 3.0 ) ( 0.0125 3.0 ) ( 0.0225 3.405 ) ( 22.5 408.0 ) ) ;

END mcon

LAYER met1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH 0.34 ;
    OFFSET 0.17 ;

    WIDTH    0.140 ;                    # Met1 1
    #SPACING  0.140 ;                    # Met1 2
    #SPACING  0.280 RANGE 3.001 100 ;	# Met1 3b
    SPACINGTABLE
	  PARALLELRUNLENGTH 0.000
	    WIDTH 0.000 0.140000
	    WIDTH 3.000000 0.280000
	    ;
    AREA 0.083 ;                        # Met1 6
    THICKNESS 0.35 ; 

    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0.000000 400.000000 ) ( 0.012500 400.000000 ) ( 0.022500 2609.000000 ) ( 22.500000 11600.000000 ) ) ;

    EDGECAPACITANCE 1.79E-6 ;
    CAPACITANCE CPERSQDIST 25.8E-6 ;
    DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
    ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
    MAXIMUMDENSITY 70.0 ;
    DENSITYCHECKWINDOW 700.0 700.0 ;
    DENSITYCHECKSTEP 70.0 ;

    RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH   0.15 ;		# Via 1a
  SPACING 0.17  ;		# Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5
  ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 ) ( 0.0125 6.0 ) ( 0.0225 6.81 ) ( 22.5 816.0 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH  0.46 ;
    OFFSET 0.23 ;

    WIDTH    0.140 ;                    # Met2 1
    #SPACING  0.140 ;                    # Met2 2
    #SPACING  0.280 RANGE 3.001 100 ;	# Met2 3b
    SPACINGTABLE
	  PARALLELRUNLENGTH 0.000
	    WIDTH 0.000 0.140000
	    WIDTH 3.000000 0.28000 ;
    AREA 0.0676 ;                       # Met2 6
    THICKNESS 0.35 ; 

    ANTENNAMODEL OXIDE1 ;
    CAPACITANCE CPERSQDIST 17.5E-6 ;
    DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
    ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 ) ( 0.0125 400.0 ) ( 0.0225 2609.0 ) ( 22.5 11600.0 ) ) ;
    
    MAXIMUMDENSITY 70.0 ;
    DENSITYCHECKWINDOW 700.0 700.0 ;
    DENSITYCHECKSTEP 70.0 ;
    RESISTANCE RPERSQ 0.125 ;
END met2

LAYER via2
  TYPE CUT ;
  WIDTH   0.20 ;		# Via2 1
  SPACING 0.20 ;		# Via2 2
  ENCLOSURE BELOW 0.040 0.085 ;	# Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ;	# Met3 4
  ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 ) ( 0.0125 6.0 ) ( 0.0225 6.81 ) ( 22.5 816.0 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC

END via2

LAYER met3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH  0.68 ;
    OFFSET 0.34 ;

    WIDTH    0.300 ;            # Met3 1
    #SPACING  0.300 ;		# Met3 2
    SPACINGTABLE
	    PARALLELRUNLENGTH 0
	    WIDTH 0 0.30
	    WIDTH 3.0 0.40 ;
    AREA     0.240 ;            # Met3 6
    THICKNESS 0.8 ;

    EDGECAPACITANCE 1.86E-6 ;
    CAPACITANCE CPERSQDIST 12.6E-6 ;
    DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
    ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 ) ( 0.0125 400.0 ) ( 0.0225 2609.0 ) ( 22.5 11600.0 ) ) ;

    MAXIMUMDENSITY 70.0 ;
    DENSITYCHECKWINDOW 700.0 700.0 ;
    DENSITYCHECKSTEP 70.0 ;
    RESISTANCE RPERSQ 0.047 ;
END met3

LAYER via3
  TYPE CUT ;

  WIDTH   0.20 ;		# Via3 1
  SPACING 0.20 ;		# Via3 2
  ENCLOSURE BELOW 0.060 0.090 ;	# Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ;	# Met4 3
  ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 ) ( 0.0125 6.0 ) ( 0.0225 6.81 ) ( 22.5 816.0 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH  0.92 ;
    OFFSET 0.46 ;

    WIDTH    0.300 ;            # Met4 1
    #SPACING  0.300 ;		# Met4 2
    
    SPACINGTABLE
	    PARALLELRUNLENGTH 0
	    WIDTH 0 0.30
	    WIDTH 3.0 0.40 ;
    AREA     0.240 ;            # Met4 4a

    THICKNESS 0.8 ;

    EDGECAPACITANCE 1.29E-6 ;
    CAPACITANCE CPERSQDIST 8.67E-6 ;
    DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
    ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 ) ( 0.0125 400.0 ) ( 0.0225 2609.0 ) ( 22.5 11600.0 ) ) ;

    MAXIMUMDENSITY 70.0 ;
    DENSITYCHECKWINDOW 700.0 700.0 ;
    DENSITYCHECKSTEP 70.0 ;
    RESISTANCE RPERSQ 0.047 ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH   0.80 ;		# Via4 1
  SPACING 0.80 ;		# Via4 2
  ENCLOSURE BELOW 0.190 0.190 ;	# Via4 4
  ENCLOSURE ABOVE 0.310 0.310 ;	# Met5 3
  ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 ) ( 0.0125 6.0 ) ( 0.0225 6.81 ) ( 22.5 816.0 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH  3.4 ;
    OFFSET 1.7 ; 

    WIDTH    1.600 ;       # Met5 1
    #SPACING  1.600 ;       # Met5 2
    SPACINGTABLE
	    PARALLELRUNLENGTH 0
	    WIDTH 0 1.600 ;
    AREA     4.000 ;       # Met5 4

    THICKNESS 1.2 ;

    ANTENNAMODEL OXIDE1 ;
    EDGECAPACITANCE 4.96E-6 ;
    CAPACITANCE CPERSQDIST 6.48E-6 ;
    DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
    ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 ) ( 0.0125 400.0 ) ( 0.0225 2609.0 ) ( 22.5 11600.0 ) ) ;
    
    RESISTANCE RPERSQ 0.0285 ;
END met5

### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER li1 ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER met1 ;
  RECT -0.145000 -0.115000 0.145000 0.115000 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0.000000 0.000000 ;
  LAYER met1 ;
  ENCLOSURE 0.060000 0.030000 ;
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  SPACING 0.360000 BY 0.360000 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER li1 ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER met1 ;
  RECT -0.115000 -0.145000 0.115000 0.145000 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0.000000 0.000000 ;
  LAYER met1 ;
  ENCLOSURE 0.030000 0.060000 ;
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  SPACING 0.360000 BY 0.360000 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER li1 ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER met1 ;
  RECT -0.115000 -0.145000 0.115000 0.145000 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0.000000 0.000000 ;
  LAYER met1 ;
  ENCLOSURE 0.030000 0.060000 ;
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  SPACING 0.360000 BY 0.360000 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER li1 ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER met1 ;
  RECT -0.145000 -0.115000 0.145000 0.115000 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0.000000 0.000000 ;
  LAYER met1 ;
  ENCLOSURE 0.060000 0.030000 ;
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  SPACING 0.360000 BY 0.360000 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER li1 ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  LAYER met1 ;
  RECT -0.145000 -0.145000 0.145000 0.145000 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0.000000 0.000000 ;
  LAYER met1 ;
  ENCLOSURE 0.060000 0.060000 ;
  LAYER mcon ;
  RECT -0.085000 -0.085000 0.085000 0.085000 ;
  SPACING 0.360000 BY 0.360000 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  LAYER met1 ;
  RECT -0.160000 -0.130000 0.160000 0.130000 ;
  LAYER met2 ;
  RECT -0.130000 -0.160000 0.130000 0.160000 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085000 0.055000 ;
  LAYER met2 ;
  ENCLOSURE 0.055000 0.085000 ;
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  SPACING 0.320000 BY 0.320000 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  LAYER met1 ;
  RECT -0.130000 -0.160000 0.130000 0.160000 ;
  LAYER met2 ;
  RECT -0.160000 -0.130000 0.160000 0.130000 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055000 0.085000 ;
  LAYER met2 ;
  ENCLOSURE 0.085000 0.055000 ;
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  SPACING 0.320000 BY 0.320000 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  LAYER met1 ;
  RECT -0.160000 -0.130000 0.160000 0.130000 ;
  LAYER met2 ;
  RECT -0.160000 -0.130000 0.160000 0.130000 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085000 0.055000 ;
  LAYER met2 ;
  ENCLOSURE 0.085000 0.055000 ;
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  SPACING 0.320000 BY 0.320000 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  LAYER met1 ;
  RECT -0.130000 -0.160000 0.130000 0.160000 ;
  LAYER met2 ;
  RECT -0.130000 -0.160000 0.130000 0.160000 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055000 0.085000 ;
  LAYER met2 ;
  ENCLOSURE 0.055000 0.085000 ;
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  SPACING 0.320000 BY 0.320000 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  LAYER met1 ;
  RECT -0.160000 -0.160000 0.160000 0.160000 ;
  LAYER met2 ;
  RECT -0.160000 -0.160000 0.160000 0.160000 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085000 0.085000 ;
  LAYER met2 ;
  ENCLOSURE 0.085000 0.085000 ;
  LAYER via ;
  RECT -0.075000 -0.075000 0.075000 0.075000 ;
  SPACING 0.320000 BY 0.320000 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met2 ;
  RECT -0.140000 -0.185000 0.140000 0.185000 ;
  LAYER met3 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.040000 0.085000 ;
  LAYER met3 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met2 ;
  RECT -0.185000 -0.140000 0.185000 0.140000 ;
  LAYER met3 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085000 0.040000 ;
  LAYER met3 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met2 ;
  RECT -0.140000 -0.185000 0.140000 0.185000 ;
  LAYER met3 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.040000 0.085000 ;
  LAYER met3 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met2 ;
  RECT -0.185000 -0.140000 0.185000 0.140000 ;
  LAYER met3 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085000 0.040000 ;
  LAYER met3 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met2 ;
  RECT -0.185000 -0.185000 0.185000 0.185000 ;
  LAYER met3 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085000 0.085000 ;
  LAYER met3 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met3 ;
  RECT -0.190000 -0.160000 0.190000 0.160000 ;
  LAYER met4 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.090000 0.060000 ;
  LAYER met4 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met3 ;
  RECT -0.160000 -0.190000 0.160000 0.190000 ;
  LAYER met4 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.060000 0.090000 ;
  LAYER met4 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met3 ;
  RECT -0.190000 -0.160000 0.190000 0.160000 ;
  LAYER met4 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.090000 0.060000 ;
  LAYER met4 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met3 ;
  RECT -0.160000 -0.190000 0.160000 0.190000 ;
  LAYER met4 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.060000 0.090000 ;
  LAYER met4 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met3 ;
  RECT -0.190000 -0.190000 0.190000 0.190000 ;
  LAYER met4 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.090000 0.090000 ;
  LAYER met4 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR_C
###  end of single via cells   ###

END LIBRARY
