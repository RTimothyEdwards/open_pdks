magic
tech sky130A
magscale 1 2
timestamp 1586352185
<< metal4 >>
rect 0 34750 200 39593
rect 0 13600 200 18593
rect 0 12410 200 13300
rect 0 11240 200 12130
rect 0 10874 200 10940
rect 0 10218 200 10814
rect 0 9922 200 10158
rect 0 9266 200 9862
rect 0 9140 200 9206
rect 0 7910 200 8840
rect 0 6940 200 7630
rect 0 5970 200 6660
rect 0 4760 200 5690
rect 0 3550 200 4480
rect 0 2580 200 3270
rect 0 1370 200 2300
rect 0 0 200 1090
<< metal5 >>
rect 0 34750 200 39593
rect 0 13600 200 18590
rect 0 12430 200 13280
rect 0 11260 200 12110
rect 0 9140 200 10940
rect 0 7930 200 8820
rect 0 6960 200 7610
rect 0 5990 200 6640
rect 0 4780 200 5670
rect 0 3570 200 4460
rect 0 2600 200 3250
rect 0 1390 200 2280
rect 0 20 200 1070
<< labels >>
flabel metal4 s 0 13600 200 18593 0 FreeSans 640 0 0 0 vddio
port 7 nsew
flabel metal5 s 0 12430 200 13280 0 FreeSans 640 0 0 0 vddio_q
port 5 nsew
flabel metal4 s 0 12410 200 13300 0 FreeSans 640 0 0 0 vddio_q
port 5 nsew
flabel metal5 s 0 11260 200 12110 0 FreeSans 640 0 0 0 vssio_q
port 11 nsew
flabel metal4 s 0 11240 200 12130 0 FreeSans 640 0 0 0 vssio_q
port 11 nsew
flabel metal5 s 0 9140 200 10940 0 FreeSans 640 0 0 0 vssa
port 2 nsew
flabel metal4 s 0 10874 200 10940 0 FreeSans 640 0 0 0 vssa
port 2 nsew
flabel metal4 s 0 10218 200 10814 0 FreeSans 640 0 0 0 amuxbus_a
port 0 nsew
flabel metal4 s 0 9266 200 9862 0 FreeSans 640 0 0 0 amuxbus_b
port 1 nsew
flabel metal4 s 0 9140 200 9206 0 FreeSans 640 0 0 0 vssa
port 2 nsew
flabel metal5 s 0 7930 200 8820 0 FreeSans 640 0 0 0 vssd
port 10 nsew
flabel metal4 s 0 7910 200 8840 0 FreeSans 640 0 0 0 vssd
port 10 nsew
flabel metal5 s 0 6960 200 7610 0 FreeSans 640 0 0 0 vssa
port 2 nsew
flabel metal4 s 0 6940 200 7630 0 FreeSans 640 0 0 0 vssa
port 2 nsew
flabel metal5 s 0 5990 200 6640 0 FreeSans 640 0 0 0 vswitch
port 4 nsew
flabel metal4 s 0 5970 200 6660 0 FreeSans 640 0 0 0 vswitch
port 4 nsew
flabel metal5 s 0 4780 200 5670 0 FreeSans 640 0 0 0 vssio
port 9 nsew
flabel metal4 s 0 4760 200 5690 0 FreeSans 640 0 0 0 vssio
port 9 nsew
flabel metal5 s 0 3570 200 4460 0 FreeSans 640 0 0 0 vddio
port 7 nsew
flabel metal4 s 0 3550 200 4480 0 FreeSans 640 0 0 0 vddio
port 7 nsew
flabel metal5 s 0 2600 200 3250 0 FreeSans 640 0 0 0 vdda
port 3 nsew
flabel metal4 s 0 2580 200 3270 0 FreeSans 640 0 0 0 vdda
port 3 nsew
flabel metal5 s 0 1390 200 2280 0 FreeSans 640 0 0 0 vccd
port 8 nsew
flabel metal4 s 0 1370 200 2300 0 FreeSans 640 0 0 0 vccd
port 8 nsew
flabel metal5 s 0 20 200 1070 0 FreeSans 640 0 0 0 vcchib
port 6 nsew
flabel metal4 s 0 0 200 1090 0 FreeSans 640 0 0 0 vcchib
port 6 nsew
flabel metal5 s 0 34750 200 39593 0 FreeSans 640 0 0 0 vssio
port 9 nsew
flabel metal5 s 0 13600 200 18590 0 FreeSans 640 0 0 0 vddio
port 7 nsew
flabel metal4 s 0 9922 200 10158 0 FreeSans 640 0 0 0 vssa
port 2 nsew
<< properties >>
string LEFclass PAD SPACER
string FIXED_BBOX 0 0 200 39593
<< end >>
