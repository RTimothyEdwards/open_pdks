VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_sc_hd__decap_20_12
  CLASS CORE SPACER ;
  FOREIGN sky130_ef_sc_hd__decap_20_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.515 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 2.200 5.430 2.635 ;
        RECT 1.670 0.630 2.010 1.460 ;
        RECT 3.490 0.950 3.840 2.200 ;
        RECT 0.085 0.085 5.430 0.630 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_ef_sc_hd__decap_20_12
END LIBRARY

