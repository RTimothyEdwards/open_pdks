magic
tech sky130A
magscale 1 2
timestamp 1602981775
<< error_p >>
rect 1389 1491 1406 1610
rect 1469 1491 1486 1610
rect 1807 1527 1815 1579
rect 1851 1527 1867 1579
rect 1998 1519 2006 1581
rect 2057 1519 2073 1581
rect 2487 1476 2523 1606
rect 2567 1476 2603 1606
rect 1878 525 1886 577
rect 1922 525 1938 577
rect 1443 486 1448 511
rect 2425 491 2429 516
rect 2732 492 2740 554
rect 2791 492 2807 554
rect 3471 538 3479 590
rect 3515 538 3531 590
<< nwell >>
rect 1134 1328 1911 1772
rect 1151 348 1976 792
rect 3212 348 3748 792
<< ndiff >>
rect 3723 1631 3986 1742
rect 2290 1476 2523 1606
rect 2567 1476 2800 1606
rect 3723 1565 3818 1631
rect 3879 1565 3986 1631
rect 3161 1510 3191 1540
rect 3723 1465 3986 1565
rect 2233 516 2404 635
rect 3816 446 3943 692
<< pdiff >>
rect 1234 1491 1406 1610
rect 1469 1491 1646 1610
rect 1251 511 1423 630
rect 3585 443 3712 689
<< psubdiff >>
rect 1998 1581 2065 1648
rect 1998 1456 2065 1519
rect 2523 1476 2567 1606
rect 2404 516 2568 635
rect 2425 453 2568 516
rect 2732 554 2799 621
rect 2732 429 2799 492
rect 3053 451 3186 695
<< nsubdiff >>
rect 1406 1491 1469 1610
rect 1807 1579 1859 1619
rect 1807 1483 1859 1527
rect 1423 511 1583 630
rect 1443 419 1583 511
rect 1878 577 1930 617
rect 1878 481 1930 525
rect 3248 446 3381 690
rect 3471 590 3523 630
rect 3471 494 3523 538
<< psubdiffcont >>
rect 1998 1519 2065 1581
rect 2732 492 2799 554
<< nsubdiffcont >>
rect 1807 1527 1859 1579
rect 1878 525 1930 577
rect 3471 538 3523 590
<< locali >>
rect 1807 1579 1859 1619
rect 1807 1483 1859 1527
rect 1998 1581 2065 1648
rect 1998 1456 2065 1519
rect 1878 577 1930 617
rect 1878 481 1930 525
rect 2732 554 2799 621
rect 3471 590 3523 630
rect 3471 494 3523 538
rect 2732 429 2799 492
<< labels >>
flabel comment s -23 575 -17 575 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s 1626 2208 1626 2208 0 FreeSans 560 0 0 0 Use_cif_see_NPLUS
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 N+_Implant_(nsd)
flabel comment s 1428 1158 1428 1158 0 FreeSans 560 0 0 0 nsd.1
flabel comment s 2568 1235 2568 1235 0 FreeSans 560 0 0 0 nsd.2
flabel comment s 1506 221 1506 221 0 FreeSans 560 0 0 0 nsd.5b
flabel comment s 2405 266 2405 266 0 FreeSans 560 0 0 0 nsd.5a
flabel comment s -39 354 -39 354 0 FreeSans 560 0 0 0 nsd.3
flabel comment s -19 185 -19 185 0 FreeSans 560 0 0 0 nsd.6
flabel comment s 3560 266 3560 266 0 FreeSans 560 0 0 0 nsd.7
flabel comment s 3291 1779 3297 1779 0 FreeSans 560 0 0 0 Incorrect
flabel comment s 3245 1364 3245 1364 0 FreeSans 560 0 0 0 nsd.10a
flabel comment s 3862 1342 3862 1342 0 FreeSans 560 0 0 0 nsd.11
flabel comment s -11 -81 -11 -81 0 FreeSans 560 0 0 0 nsd.9
flabel comment s 15 48 15 48 0 FreeSans 560 0 0 0 nsd.8
<< end >>
