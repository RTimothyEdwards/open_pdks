magic
tech s8seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
tri 530 2319 590 2344 se
tri 590 2319 615 2344 sw
tri 530 2234 615 2319 ne
tri 615 2234 700 2319 sw
tri 615 2149 700 2234 ne
tri 700 2149 785 2234 sw
tri 700 2064 785 2149 ne
tri 785 2064 870 2149 sw
tri 785 1979 870 2064 ne
tri 870 1979 955 2064 sw
tri 870 1894 955 1979 ne
tri 955 1894 1040 1979 sw
tri 955 1809 1040 1894 ne
tri 1040 1809 1125 1894 sw
tri 1040 1724 1125 1809 ne
tri 1125 1724 1210 1809 sw
tri 1125 1639 1210 1724 ne
tri 1210 1639 1295 1724 sw
tri 1210 1554 1295 1639 ne
tri 1295 1554 1380 1639 sw
tri 1295 1469 1380 1554 ne
tri 1380 1469 1465 1554 sw
tri 1380 1384 1465 1469 ne
tri 1465 1384 1550 1469 sw
tri 1465 1299 1550 1384 ne
tri 1550 1299 1635 1384 sw
tri 1550 1214 1635 1299 ne
tri 1635 1214 1720 1299 sw
tri 1635 1129 1720 1214 ne
tri 1720 1129 1805 1214 sw
tri 1720 1044 1805 1129 ne
tri 1805 1044 1890 1129 sw
tri 1805 959 1890 1044 ne
tri 1890 959 1975 1044 sw
tri 1890 874 1975 959 ne
tri 1975 874 2060 959 sw
tri 1975 789 2060 874 ne
tri 2060 789 2145 874 sw
tri 2060 704 2145 789 ne
tri 2145 704 2230 789 sw
tri 2145 619 2230 704 ne
tri 2230 619 2315 704 sw
tri 2230 534 2315 619 ne
tri 2315 590 2344 619 sw
rect 2315 534 51200 590
tri 2315 530 2319 534 ne
rect 2319 530 51200 534
<< end >>
