
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;

SITE unit
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE  0.480 BY 3.400 ;
END unit

######  Starting overlap layers #####
# ******** Layer OverlapCheck, type blockage, number 90 **************
LAYER OverlapCheck
  TYPE OVERLAP ;
END OverlapCheck

######  Starting routing layers - metal and via #####
# ******** Layer li1, type routing, number 56 **************
LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.48 ;
  MINWIDTH 0.170000 ;
  WIDTH 0.170000 ;
  AREA 0.028900 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0 0.170000 ;
  THICKNESS 0.100000 ;
  EDGECAPACITANCE 3.26E-6 ;
  CAPACITANCE CPERSQDIST 36.9E-6 ;
  RESISTANCE RPERSQ 12.2 ;
#  DCCURRENTDENSITY AVERAGE (no limit on this layer) ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0.000000 75.000000 ) ( 0.012500 75.000000 ) ( 0.022500 85.125000 ) ( 22.500000 10200.000000 ) ) ;
END li1

# ******** Layer mcon, type routing, number 35 **************
LAYER mcon
  TYPE CUT ;
  SPACING 0.190000 ;
  WIDTH 0.170000 ;
  ANTENNADIFFAREARATIO PWL ( ( 0.000000 3.000000 ) ( 0.012500 3.000000 ) ( 0.022500 3.405000 ) ( 22.500000 408.000000 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC
  ENCLOSURE BELOW 0.000000 0.000000 ;
  ENCLOSURE ABOVE 0.000000 0.000000 ;
END mcon

# ******** Layer met1, type routing, number 36 **************
LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.37 ;
  MINENCLOSEDAREA 0.140000 ;
  MINWIDTH 0.140000 ;
  WIDTH 0.140000 ;
  AREA 0.083000 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.000
    WIDTH 0.000 0.140000
    WIDTH 3.000000 0.280000
    ;
  THICKNESS 0.350000 ;
  EDGECAPACITANCE 1.79E-6 ;
  CAPACITANCE CPERSQDIST 25.8E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0.000000 400.000000 ) ( 0.012500 400.000000 ) ( 0.022500 2609.000000 ) ( 22.500000 11600.000000 ) ) ;
END met1

# ******** Layer via, type routing, number 40 **************
LAYER via1
  TYPE CUT ;
  SPACING 0.170000 ;
  WIDTH 0.150000 ;
  ANTENNADIFFAREARATIO PWL ( ( 0.000000 6.000000 ) ( 0.012500 6.000000 ) ( 0.022500 6.810000 ) ( 22.500000 816.000000 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
  ENCLOSURE BELOW 0.000000 0.000000 ;
  ENCLOSURE ABOVE 0.000000 0.000000 ;
END via1

# ******** Layer met2, type routing, number 41 **************
LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.48 ;
  MINENCLOSEDAREA 0.140000 ;
  MINWIDTH 0.140000 ;
  WIDTH 0.140000 ;
  AREA 0.067600 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.000
    WIDTH 0.000 0.140000
    WIDTH 3.000000 0.280000
    ;
  THICKNESS 0.350000 ;
  EDGECAPACITANCE 1.22E-6 ;
  CAPACITANCE CPERSQDIST 17.5E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0.000000 400.000000 ) ( 0.012500 400.000000 ) ( 0.022500 2609.000000 ) ( 22.500000 11600.000000 ) ) ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  SPACING 0.200000 ;
  WIDTH 0.200000 ;
  ANTENNADIFFAREARATIO PWL ( ( 0.000000 6.000000 ) ( 0.012500 6.000000 ) ( 0.022500 6.810000 ) ( 22.500000 816.000000 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
  ENCLOSURE BELOW 0.000000 0.000000 ;
  ENCLOSURE ABOVE 0.000000 0.000000 ;
END via2

# ******** Layer met3, type routing, number 34 **************
LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.666 ;
  MINWIDTH 0.300000 ;
  WIDTH 0.300000 ;
  AREA 0.240000 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.000
    WIDTH 0.000 0.300000
    WIDTH 3.000000 0.400000
    ;
  THICKNESS 0.800000 ;
  EDGECAPACITANCE 1.86E-6 ;
  CAPACITANCE CPERSQDIST 12.6E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0.000000 400.000000 ) ( 0.012500 400.000000 ) ( 0.022500 2609.000000 ) ( 22.500000 11600.000000 ) ) ;
END met3

# ******** Layer via3, type routing, number 70 **************
LAYER via3
  TYPE CUT ;
  SPACING 0.200000 ;
  WIDTH 0.200000 ;
  ANTENNADIFFAREARATIO PWL ( ( 0.000000 6.000000 ) ( 0.012500 6.000000 ) ( 0.022500 6.810000 ) ( 22.500000 816.000000 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
  ENCLOSURE BELOW 0.000000 0.000000 ;
  ENCLOSURE ABOVE 0.000000 0.000000 ;
END via3

# ******** Layer met4, type routing, number 71 **************
LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.96 ;
  MINWIDTH 0.300000 ;
  WIDTH 0.300000 ;
  AREA 0.240000 ;
  SPACINGTABLE
  PARALLELRUNLENGTH 0.000
    WIDTH 0.000 0.300000
    WIDTH 3.000000 0.400000
    ;
  THICKNESS 0.800000 ;
  EDGECAPACITANCE 1.29E-6 ;
  CAPACITANCE CPERSQDIST 8.67E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0.000000 400.000000 ) ( 0.012500 400.000000 ) ( 0.022500 2609.000000 ) ( 22.500000 11600.000000 ) ) ;
END met4

# ******** Layer via4, type routing, number 58 **************
LAYER via4
  TYPE CUT ;
  SPACING 0.800000 ;
  WIDTH 0.800000 ;
  ANTENNADIFFAREARATIO PWL ( ( 0.000000 6.000000 ) ( 0.012500 6.000000 ) ( 0.022500 6.810000 ) ( 22.500000 816.000000 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
  ENCLOSURE BELOW 0.000000 0.000000 ;
  ENCLOSURE ABOVE 0.000000 0.000000 ;
END via4

# ******** Layer met5, type routing, number 72 **************
LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.3 ;
  MINWIDTH 1.600000 ;
  WIDTH 1.600000 ;
  AREA 2.560000 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0
    WIDTH 0 1.600000 ;
  THICKNESS 1.200000 ;
  EDGECAPACITANCE 4.96E-6 ;
  CAPACITANCE CPERSQDIST 6.48E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0.000000 400.000000 ) ( 0.012500 400.000000 ) ( 0.022500 2609.000000 ) ( 22.500000 11600.000000 ) ) ;
END met5

######  completed routing layers - metal and via #####

### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 LAYER li1 ;
 RECT -0.085 -0.165 0.085 0.165 ;
 LAYER met1 ;
 RECT -0.16 -0.13 0.16 0.13 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
 LAYER li1 ;
 ENCLOSURE 0.000 0.080 ;
 LAYER met1 ;
 ENCLOSURE 0.030 0.060 ;
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 SPACING 0.360 BY 0.360 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 LAYER li1 ;
 RECT -0.165 -0.085 0.165 0.085 ;
 LAYER met1 ;
 RECT -0.13 -0.16 0.13 0.16 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
 LAYER li1 ;
 ENCLOSURE 0.000 0.080 ;
 LAYER met1 ;
 ENCLOSURE 0.030 0.060 ;
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 SPACING 0.360 BY 0.360 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 LAYER li1 ;
 RECT -0.085 -0.165 0.085 0.165 ;
 LAYER met1 ;
 RECT -0.13 -0.16 0.13 0.16 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
 LAYER li1 ;
 ENCLOSURE 0.000 0.080 ;
 LAYER met1 ;
 ENCLOSURE 0.030 0.060 ;
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 SPACING 0.360 BY 0.360 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 LAYER li1 ;
 RECT -0.165 -0.085 0.165 0.085 ;
 LAYER met1 ;
 RECT -0.16 -0.13 0.16 0.13 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
 LAYER li1 ;
 ENCLOSURE 0.000 0.080 ;
 LAYER met1 ;
 ENCLOSURE 0.030 0.060 ;
 LAYER mcon ;
 RECT -0.085 -0.085 0.085 0.085 ;
 SPACING 0.360 BY 0.360 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
# VIA L1M1_PR_C DEFAULT
#   LAYER mcon ;
#   RECT -0.085000 -0.085000 0.085000 0.085000 ;
#   LAYER li1 ;
#   RECT -0.085000 -0.085000 0.085000 0.085000 ;
#   LAYER met1 ;
#   RECT -0.145000 -0.145000 0.145000 0.145000 ;
# END L1M1_PR_C

# VIARULE L1M1_PR_C GENERATE
#   LAYER li1 ;
#   ENCLOSURE 0.000000 0.000000 ;
#   LAYER met1 ;
#   ENCLOSURE 0.060000 0.060000 ;
#   LAYER mcon ;
#   RECT -0.085000 -0.085000 0.085000 0.085000 ;
#   SPACING 0.360000 BY 0.360000 ;
# END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 LAYER met1 ;
 RECT -0.16 -0.13 0.16 0.13 ;
 LAYER met2 ;
 RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
 LAYER met1 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER met2 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 SPACING 0.320 BY 0.320 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 LAYER met1 ;
 RECT -0.13 -0.16 0.13 0.16 ;
 LAYER met2 ;
 RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
 LAYER met1 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER met2 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 SPACING 0.320 BY 0.320 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 LAYER met1 ;
 RECT -0.16 -0.13 0.16 0.13 ;
 LAYER met2 ;
 RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
 LAYER met1 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER met2 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 SPACING 0.320 BY 0.320 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 LAYER met1 ;
 RECT -0.13 -0.16 0.13 0.16 ;
 LAYER met2 ;
 RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
 LAYER met1 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER met2 ;
 ENCLOSURE 0.055 0.085 ;
 LAYER via1 ;
 RECT -0.075 -0.075 0.075 0.075 ;
 SPACING 0.320 BY 0.320 ;
END M1M2_PR_MR

# # Centered via rule, we really do not want to use it
# VIA M1M2_PR_C DEFAULT
#   LAYER via ;
#   RECT -0.075000 -0.075000 0.075000 0.075000 ;
#   LAYER met1 ;
#   RECT -0.160000 -0.160000 0.160000 0.160000 ;
#   LAYER met2 ;
#   RECT -0.160000 -0.160000 0.160000 0.160000 ;
# END M1M2_PR_C

# VIARULE M1M2_PR_C GENERATE
#   LAYER met1 ;
#   ENCLOSURE 0.085000 0.085000 ;
#   LAYER met2 ;
#   ENCLOSURE 0.085000 0.085000 ;
#   LAYER via ;
#   RECT -0.075000 -0.075000 0.075000 0.075000 ;
#   SPACING 0.320000 BY 0.320000 ;
# END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
 LAYER via2 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 LAYER met2 ;
 RECT -0.14 -0.185 0.14 0.185 ;
 LAYER met3 ;
 RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
 LAYER met2 ;
 ENCLOSURE 0.040 0.085 ;
 LAYER met3 ;
 ENCLOSURE 0.065 0.065 ;
 LAYER via2 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 SPACING 0.40 BY 0.40 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
 LAYER via2 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 LAYER met2 ;
 RECT -0.185 -0.14 0.185 0.14 ;
 LAYER met3 ;
 RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
 LAYER met2 ;
 ENCLOSURE 0.040 0.085 ;
 LAYER met3 ;
 ENCLOSURE 0.065 0.065 ;
 LAYER via2 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 SPACING 0.40 BY 0.40 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met2 ;
  RECT -0.140000 -0.185000 0.140000 0.185000 ;
  LAYER met3 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.040000 0.085000 ;
  LAYER met3 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met2 ;
  RECT -0.185000 -0.140000 0.185000 0.140000 ;
  LAYER met3 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085000 0.040000 ;
  LAYER met3 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via2 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M2M3_PR_MR

# # Centered via rule, we really do not want to use it
# VIA M2M3_PR_C DEFAULT
#   LAYER via2 ;
#   RECT -0.100000 -0.100000 0.100000 0.100000 ;
#   LAYER met2 ;
#   RECT -0.185000 -0.185000 0.185000 0.185000 ;
#   LAYER met3 ;
#   RECT -0.165000 -0.165000 0.165000 0.165000 ;
# END M2M3_PR_C

# VIARULE M2M3_PR_C GENERATE
#   LAYER met2 ;
#   ENCLOSURE 0.085000 0.085000 ;
#   LAYER met3 ;
#   ENCLOSURE 0.065000 0.065000 ;
#   LAYER via2 ;
#   RECT -0.100000 -0.100000 0.100000 0.100000 ;
#   SPACING 0.400000 BY 0.400000 ;
# END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
 LAYER via3 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 LAYER met3 ;
 RECT -0.19 -0.16 0.19 0.16 ;
 LAYER met4 ;
 RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
 LAYER met3 ;
 ENCLOSURE 0.06 0.09 ;
 LAYER met4 ;
 ENCLOSURE 0.065 0.065 ;
 LAYER via3 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 SPACING 0.40 BY 0.40 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
 LAYER via3 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 LAYER met3 ;
 RECT -0.16 -0.19 0.16 0.19 ;
 LAYER met4 ;
 RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
 LAYER met3 ;
 ENCLOSURE 0.06 0.09 ;
 LAYER met4 ;
 ENCLOSURE 0.065 0.065 ;
 LAYER via3 ;
 RECT -0.1 -0.1 0.1 0.1 ;
 SPACING 0.40 BY 0.40 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met3 ;
  RECT -0.190000 -0.160000 0.190000 0.160000 ;
  LAYER met4 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.090000 0.060000 ;
  LAYER met4 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  LAYER met3 ;
  RECT -0.160000 -0.190000 0.160000 0.190000 ;
  LAYER met4 ;
  RECT -0.165000 -0.165000 0.165000 0.165000 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.060000 0.090000 ;
  LAYER met4 ;
  ENCLOSURE 0.065000 0.065000 ;
  LAYER via3 ;
  RECT -0.100000 -0.100000 0.100000 0.100000 ;
  SPACING 0.400000 BY 0.400000 ;
END M3M4_PR_MR

# # Centered via rule, we really do not want to use it
# VIA M3M4_PR_C DEFAULT
#   LAYER via3 ;
#   RECT -0.100000 -0.100000 0.100000 0.100000 ;
#   LAYER met3 ;
#   RECT -0.190000 -0.190000 0.190000 0.190000 ;
#   LAYER met4 ;
#   RECT -0.165000 -0.165000 0.165000 0.165000 ;
# END M3M4_PR_C

# VIARULE M3M4_PR_C GENERATE
#   LAYER met3 ;
#   ENCLOSURE 0.090000 0.090000 ;
#   LAYER met4 ;
#   ENCLOSURE 0.065000 0.065000 ;
#   LAYER via3 ;
#   RECT -0.100000 -0.100000 0.100000 0.100000 ;
#   SPACING 0.400000 BY 0.400000 ;
# END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
 LAYER via4 ;
 RECT -0.4 -0.4 0.4 0.4 ;
 LAYER met4 ;
 RECT -0.59 -0.59 0.59 0.59 ;
 LAYER met5 ;
 RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
 LAYER met4 ;
 ENCLOSURE 0.190 0.190 ;
 LAYER met5 ;
 ENCLOSURE 0.310 0.310 ;
 LAYER via4 ;
 RECT -0.4 -0.4 0.4 0.4 ;
 SPACING 1.60 BY 1.60 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER met4 ;
  RECT -0.590000 -0.590000 0.590000 0.590000 ;
  LAYER met5 ;
  RECT -0.710000 -0.710000 0.710000 0.710000 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.190000 0.190000 ;
  LAYER met5 ;
  ENCLOSURE 0.310000 0.310000 ;
  LAYER via4 ;
  RECT -0.400000 -0.400000 0.400000 0.400000 ;
  SPACING 1.600000 BY 1.600000 ;
END M4M5_PR_MR

# # Centered via rule, we really do not want to use it
# VIA M4M5_PR_C DEFAULT
#   LAYER via4 ;
#   RECT -0.400000 -0.400000 0.400000 0.400000 ;
#   LAYER met4 ;
#   RECT -0.590000 -0.590000 0.590000 0.590000 ;
#   LAYER met5 ;
#   RECT -0.710000 -0.710000 0.710000 0.710000 ;
# END M4M5_PR_C

# VIARULE M4M5_PR_C GENERATE
#   LAYER met4 ;
#   ENCLOSURE 0.190000 0.190000 ;
#   LAYER met5 ;
#   ENCLOSURE 0.310000 0.310000 ;
#   LAYER via4 ;
#   RECT -0.400000 -0.400000 0.400000 0.400000 ;
#   SPACING 1.600000 BY 1.600000 ;
# END M4M5_PR_C

END LIBRARY
