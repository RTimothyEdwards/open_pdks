magic
tech sky130A
magscale 1 2
timestamp 1602981889
<< error_p >>
rect 3687 1776 4022 1778
rect 3723 1740 3986 1742
rect 1389 1491 1406 1610
rect 1469 1491 1486 1610
rect 1807 1527 1815 1579
rect 1851 1527 1867 1579
rect 1998 1519 2006 1581
rect 2057 1519 2073 1581
rect 2487 1476 2523 1606
rect 2567 1476 2603 1606
rect 1878 525 1886 577
rect 1922 525 1938 577
rect 1438 486 1448 511
rect 2420 491 2429 516
rect 2732 492 2740 554
rect 2791 492 2807 554
rect 3441 538 3449 590
rect 3485 538 3501 590
<< nwell >>
rect 1922 1322 4125 1776
rect 2098 348 3210 792
rect 3750 350 4194 794
<< ndiff >>
rect 1234 1491 1406 1610
rect 1469 1491 1646 1610
rect 1251 511 1423 630
rect 3555 443 3682 689
<< pdiff >>
rect 3723 1631 3986 1742
rect 2290 1476 2523 1606
rect 2567 1476 2800 1606
rect 3723 1565 3818 1631
rect 3879 1565 3986 1631
rect 3161 1510 3191 1540
rect 3723 1465 3986 1565
rect 2233 516 2404 635
rect 3786 446 3913 692
<< psubdiff >>
rect 1406 1491 1469 1610
rect 1807 1579 1859 1619
rect 1807 1483 1859 1527
rect 1423 511 1578 630
rect 1438 419 1578 511
rect 1878 577 1930 617
rect 1878 481 1930 525
rect 3236 446 3369 690
rect 3441 590 3493 630
rect 3441 494 3493 538
<< nsubdiff >>
rect 1998 1581 2065 1648
rect 1998 1456 2065 1519
rect 2523 1476 2567 1606
rect 2404 516 2563 635
rect 2420 453 2563 516
rect 2732 554 2799 621
rect 2732 429 2799 492
rect 3041 451 3174 695
<< psubdiffcont >>
rect 1807 1527 1859 1579
rect 1878 525 1930 577
rect 3441 538 3493 590
<< nsubdiffcont >>
rect 1998 1519 2065 1581
rect 2732 492 2799 554
<< locali >>
rect 1807 1579 1859 1619
rect 1807 1483 1859 1527
rect 1998 1581 2065 1648
rect 1998 1456 2065 1519
rect 1878 577 1930 617
rect 1878 481 1930 525
rect 2732 554 2799 621
rect 3441 590 3493 630
rect 3441 494 3493 538
rect 2732 429 2799 492
<< labels >>
flabel comment s 3291 1779 3297 1779 0 FreeSans 560 0 0 0 Incorrect
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 P+_Implant_(psd)
flabel comment s 1428 1158 1428 1158 0 FreeSans 560 0 0 0 psd.1
flabel comment s 2568 1235 2568 1235 0 FreeSans 560 0 0 0 psd.2
flabel comment s 3245 1364 3245 1364 0 FreeSans 560 0 0 0 psd.10a
flabel comment s 3862 1342 3862 1342 0 FreeSans 560 0 0 0 psd.11
flabel comment s 1506 221 1506 221 0 FreeSans 560 0 0 0 psd.5b
flabel comment s 2405 266 2405 266 0 FreeSans 560 0 0 0 psd.5a
flabel comment s 3560 266 3560 266 0 FreeSans 560 0 0 0 psd.7
flabel comment s 1626 2208 1626 2208 0 FreeSans 560 0 0 0 Use_cif_see_PPLUS
flabel comment s 165 1261 171 1261 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s 169 871 169 871 0 FreeSans 560 0 0 0 psd.6
flabel comment s 149 1040 149 1040 0 FreeSans 560 0 0 0 psd.3
flabel comment s 178 603 178 603 0 FreeSans 560 0 0 0 psd.9
flabel comment s 173 758 173 758 0 FreeSans 560 0 0 0 psd.8
<< end >>
