VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__top_xres4v2
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_xres4v2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY R90 ;
  PIN PAD_A_ESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.245 0.000 18.910 0.565 ;
    END
    PORT
      LAYER met2 ;
        RECT 17.245 0.000 18.910 0.565 ;
    END
  END PAD_A_ESD_H
  PIN XRES_H_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.935 0.000 29.665 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.935 0.000 29.665 0.330 ;
    END
  END XRES_H_N
  PIN FILT_IN_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.075 0.000 21.225 1.410 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.075 0.000 21.225 1.410 ;
    END
  END FILT_IN_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.400 0.000 8.920 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 8.425 0.000 8.895 0.330 ;
    END
  END ENABLE_VDDIO
  PIN TIE_WEAK_HI_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.190 0.000 73.260 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 72.215 0.000 73.235 0.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 49.985 73.925 64.465 ;
    END
  END TIE_WEAK_HI_H
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.285 0.000 12.545 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 12.285 0.000 12.545 0.330 ;
    END
  END ENABLE_H
  PIN PULLUP_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.555 0.000 15.135 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 14.555 0.000 15.135 0.330 ;
    END
  END PULLUP_H
  PIN EN_VDDIO_SIG_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.360 0.000 22.660 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.360 0.000 22.660 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320 5.360 29.580 10.980 ;
    END
  END EN_VDDIO_SIG_H
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.580 0.000 28.230 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.580 0.000 28.230 0.330 ;
    END
  END TIE_LO_ESD
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.505 0.000 31.155 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 30.505 0.000 31.155 0.330 ;
    END
  END TIE_HI_ESD
  PIN DISABLE_PULLUP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.760 0.000 33.020 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 32.760 0.000 33.020 0.330 ;
    END
  END DISABLE_PULLUP_H
  PIN INP_SEL_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.905 0.000 25.135 9.975 ;
    END
  END INP_SEL_H
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
  END VSSIO
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
  END VSSD
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
  END VDDIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
  END VSWITCH
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
  END VCCHIB
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
  END VSSIO_Q
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 17.250 108.455 54.435 164.285 ;
    END
  END PAD
  OBS
      LAYER nwell ;
        RECT -0.515 168.515 75.620 170.210 ;
        RECT -0.515 146.690 1.675 168.515 ;
        RECT 73.095 146.690 75.620 168.515 ;
        RECT -0.515 144.880 75.620 146.690 ;
      LAYER pwell ;
        RECT -0.290 140.685 75.290 144.565 ;
      LAYER nwell ;
        RECT -0.330 130.665 75.330 140.380 ;
      LAYER pwell ;
        RECT -0.130 129.315 41.750 130.355 ;
        RECT 61.910 129.315 75.130 130.355 ;
        RECT -0.130 124.135 75.130 129.315 ;
        RECT -0.130 102.525 1.435 124.135 ;
        RECT 73.560 102.525 75.130 124.135 ;
        RECT -0.130 99.230 75.130 102.525 ;
        RECT -0.130 97.995 58.470 99.230 ;
        RECT 71.930 97.995 75.130 99.230 ;
        RECT -0.130 96.735 75.130 97.995 ;
        RECT -0.130 96.730 58.470 96.735 ;
      LAYER li1 ;
        RECT 0.000 144.435 75.000 199.220 ;
        RECT -0.160 140.815 75.160 144.435 ;
        RECT 0.000 130.225 75.000 140.815 ;
        RECT -0.265 101.395 75.000 130.225 ;
        RECT 0.000 0.185 75.000 101.395 ;
      LAYER met1 ;
        RECT 0.000 170.090 75.000 199.210 ;
        RECT -0.145 131.275 75.145 170.090 ;
        RECT 0.000 130.220 75.000 131.275 ;
        RECT -0.145 95.895 75.145 130.220 ;
        RECT 0.000 10.255 75.000 95.895 ;
        RECT 0.000 0.610 24.625 10.255 ;
        RECT 0.000 0.185 12.005 0.610 ;
        RECT 12.825 0.185 14.275 0.610 ;
        RECT 15.415 0.185 22.080 0.610 ;
        RECT 22.940 0.185 24.625 0.610 ;
        RECT 25.415 0.610 75.000 10.255 ;
        RECT 25.415 0.185 27.300 0.610 ;
        RECT 28.510 0.185 30.225 0.610 ;
        RECT 31.435 0.185 32.480 0.610 ;
        RECT 33.300 0.185 75.000 0.610 ;
      LAYER met2 ;
        RECT 0.340 11.260 74.915 199.210 ;
        RECT 0.340 5.080 29.040 11.260 ;
        RECT 29.860 5.080 74.915 11.260 ;
        RECT 0.340 1.690 74.915 5.080 ;
        RECT 0.340 0.845 19.795 1.690 ;
        RECT 0.340 0.610 16.965 0.845 ;
        RECT 0.340 0.000 8.145 0.610 ;
        RECT 9.175 0.000 12.005 0.610 ;
        RECT 12.825 0.000 14.275 0.610 ;
        RECT 15.415 0.000 16.965 0.610 ;
        RECT 19.190 0.000 19.795 0.845 ;
        RECT 21.505 0.610 74.915 1.690 ;
        RECT 21.505 0.000 22.080 0.610 ;
        RECT 22.940 0.000 27.300 0.610 ;
        RECT 28.510 0.000 28.655 0.610 ;
        RECT 29.945 0.000 30.225 0.610 ;
        RECT 31.435 0.000 32.480 0.610 ;
        RECT 33.300 0.000 71.935 0.610 ;
        RECT 73.515 0.000 74.915 0.610 ;
      LAYER met3 ;
        RECT 0.965 64.865 74.700 200.000 ;
        RECT 0.965 49.585 71.790 64.865 ;
        RECT 74.325 49.585 74.700 64.865 ;
        RECT 0.965 1.810 74.700 49.585 ;
        RECT 0.965 0.965 19.675 1.810 ;
        RECT 0.965 0.730 16.845 0.965 ;
        RECT 0.965 0.330 8.000 0.730 ;
        RECT 9.320 0.330 16.845 0.730 ;
        RECT 19.310 0.330 19.675 0.965 ;
        RECT 21.625 0.730 74.700 1.810 ;
        RECT 21.625 0.330 28.535 0.730 ;
        RECT 30.065 0.330 71.790 0.730 ;
        RECT 73.660 0.330 74.700 0.730 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 165.885 75.000 174.185 ;
        RECT 0.000 106.855 15.650 165.885 ;
        RECT 56.035 106.855 75.000 165.885 ;
        RECT 0.000 96.585 75.000 106.855 ;
        RECT 2.870 18.285 72.130 96.585 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__top_xres4v2
END LIBRARY

