magic
tech s8seal_ring
magscale 1 2
timestamp 1584558827
<< type65_20 >>
rect 290 2244 350 51210
tri 290 2219 350 2244 nw
<< end >>
