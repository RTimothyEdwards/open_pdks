magic
tech s8seal_ring
magscale 1 2
timestamp 1584558827
<< type81_1 >>
rect 0 2597 1200 51210
tri 0 0 1200 2597 nw
<< end >>
