magic
tech sky130A
magscale 1 2
timestamp 1609170569
<< metal3 >>
rect 2908 38501 4894 38507
rect 2908 34872 2914 38501
rect 4888 34872 4894 38501
rect 5280 38501 7266 38507
rect 5280 34882 5286 38501
rect 7260 34882 7266 38501
rect 5280 34876 7266 34882
rect 2908 34866 4894 34872
rect 7624 18544 9746 18550
rect 7624 13650 7630 18544
rect 9740 13650 9746 18544
rect 7624 13644 9746 13650
rect 5216 5654 7336 5660
rect 5216 4798 5222 5654
rect 7330 4798 7336 5654
rect 5216 4792 7336 4798
rect 7604 4444 9750 4450
rect 7604 3590 7610 4444
rect 9744 3590 9750 4444
rect 7604 3584 9750 3590
<< via3 >>
rect 2914 34872 4888 38501
rect 5286 34882 7260 38501
rect 7630 13650 9740 18544
rect 5222 4798 7330 5654
rect 7610 3590 9744 4444
<< metal4 >>
rect 2908 34872 2914 38501
rect 4888 34872 4894 38501
rect 5280 34882 5286 38501
rect 7260 34882 7266 38501
rect 5280 34876 7266 34882
rect 2908 34866 4894 34872
rect 7624 18544 9746 18550
rect 7624 13650 7630 18544
rect 9740 13650 9746 18544
rect 7624 13644 9746 13650
rect 5216 5654 7336 5660
rect 5216 4798 5222 5654
rect 7330 4798 7336 5654
rect 5216 4792 7336 4798
rect 7604 4444 9750 4450
rect 7604 3590 7610 4444
rect 9744 3590 9750 4444
rect 7604 3584 9750 3590
<< properties >>
string FIXED_BBOX 0 -406 15000 39592
<< end >>
