magic
tech sky130A
magscale 1 2
timestamp 1584383567
<< error_s >>
rect 119603 132136 121521 132218
rect 98716 131466 98782 131482
rect 800 131078 866 131094
rect 1823 129308 1824 129332
rect 1904 129308 1905 129332
rect 2377 129308 2378 129332
rect 2458 129308 2459 129332
rect 2931 129308 2932 129332
rect 3012 129308 3013 129332
rect 3485 129308 3486 129332
rect 3566 129308 3567 129332
rect 4039 129308 4040 129332
rect 4120 129308 4121 129332
rect 4593 129308 4594 129332
rect 4674 129308 4675 129332
rect 5147 129308 5148 129332
rect 5228 129308 5229 129332
rect 5701 129308 5702 129332
rect 5782 129308 5783 129332
rect 6255 129308 6256 129332
rect 6336 129308 6337 129332
rect 6809 129308 6810 129332
rect 6890 129308 6891 129332
rect 7363 129308 7364 129332
rect 7444 129308 7445 129332
rect 7917 129308 7918 129332
rect 7998 129308 7999 129332
rect 8471 129308 8472 129332
rect 8552 129308 8553 129332
rect 9025 129308 9026 129332
rect 9106 129308 9107 129332
rect 9579 129308 9580 129332
rect 9660 129308 9661 129332
rect 10133 129308 10134 129332
rect 10214 129308 10215 129332
rect 10687 129308 10688 129332
rect 10768 129308 10769 129332
rect 11241 129308 11242 129332
rect 11322 129308 11323 129332
rect 11795 129308 11796 129332
rect 11876 129308 11877 129332
rect 12349 129308 12350 129332
rect 12430 129308 12431 129332
rect 1847 129284 1881 129296
rect 2401 129284 2435 129296
rect 2955 129284 2989 129296
rect 3509 129284 3543 129296
rect 4063 129284 4097 129296
rect 4617 129284 4651 129296
rect 5171 129284 5205 129296
rect 5725 129284 5759 129296
rect 6279 129284 6313 129296
rect 6833 129284 6867 129296
rect 7387 129284 7421 129296
rect 7941 129284 7975 129296
rect 8495 129284 8529 129296
rect 9049 129284 9083 129296
rect 9603 129284 9637 129296
rect 10157 129284 10191 129296
rect 10711 129284 10745 129296
rect 11265 129284 11299 129296
rect 11819 129284 11853 129296
rect 12373 129284 12407 129296
rect 22784 129100 22856 131100
rect 23055 129133 23173 131027
rect 23444 129100 23504 131100
rect 23704 129100 23776 131100
rect 23975 129133 24093 131027
rect 24364 129100 24424 131100
rect 24624 129100 24696 131100
rect 24895 129133 25013 131027
rect 25284 129100 25344 131100
rect 25544 129100 25616 131100
rect 25815 129133 25933 131027
rect 26204 129100 26264 131100
rect 26464 129100 26536 131100
rect 26735 129133 26853 131027
rect 27124 129100 27184 131100
rect 27384 129100 27456 131100
rect 27655 129133 27773 131027
rect 28044 129100 28104 131100
rect 28304 129100 28376 131100
rect 28575 129133 28693 131027
rect 28964 129100 29024 131100
rect 29224 129100 29296 131100
rect 29495 129133 29613 131027
rect 29884 129100 29944 131100
rect 30144 129100 30216 131100
rect 30415 129133 30533 131027
rect 30804 129100 30864 131100
rect 31064 129100 31136 131100
rect 31335 129133 31453 131027
rect 31724 129100 31784 131100
rect 31984 129100 32056 131100
rect 32255 129133 32373 131027
rect 32644 129100 32704 131100
rect 119390 131001 119472 132035
rect 119682 131171 119764 131865
rect 119904 131854 121210 131936
rect 120072 131660 121014 131710
rect 119941 131617 119967 131628
rect 119957 131577 120051 131617
rect 120963 131577 121057 131617
rect 119957 131417 120051 131457
rect 120963 131417 121057 131457
rect 119941 131406 119967 131417
rect 120072 131316 121014 131366
rect 119904 131102 121210 131184
rect 121250 131171 121332 131865
rect 121542 131001 121624 132035
rect 122443 131134 122493 132134
rect 122593 131134 122721 132134
rect 122749 131134 122799 132134
rect 122865 131134 122915 132134
rect 123075 131134 123131 132134
rect 123291 131134 123347 132134
rect 123447 131134 123575 132134
rect 123603 131134 123653 132134
rect 123769 131134 123819 132134
rect 123979 131134 124035 132134
rect 124135 131134 124263 132134
rect 124291 131134 124347 132134
rect 124447 131134 124575 132134
rect 124603 131134 124659 132134
rect 124759 131134 124809 132134
rect 124875 131134 124925 131734
rect 125025 131134 125075 131734
rect 125141 131134 125191 132134
rect 125291 131134 125347 132134
rect 125447 131134 125497 132134
rect 126387 131130 126445 131164
rect 127227 131142 127277 132142
rect 127377 131142 127505 132142
rect 127533 131142 127661 132142
rect 127689 131142 127817 132142
rect 127845 131142 127973 132142
rect 128001 131142 128051 132142
rect 128117 131142 128167 132142
rect 128267 131142 128323 132142
rect 128423 131142 128473 132142
rect 128539 131142 128589 132142
rect 128689 131142 128817 132142
rect 128845 131142 128901 132142
rect 129001 131142 129129 132142
rect 129157 131142 129207 132142
rect 129273 131142 129323 132142
rect 129423 131142 129551 132142
rect 129579 131142 129635 132142
rect 129735 131142 129863 132142
rect 129891 131514 129941 132142
rect 129891 131442 129944 131514
rect 129891 131142 129941 131442
rect 130004 131142 130016 131442
rect 133592 130979 134592 131029
rect 39774 130302 39840 130318
rect 40797 128532 40798 128556
rect 40878 128532 40879 128556
rect 41351 128532 41352 128556
rect 41432 128532 41433 128556
rect 41905 128532 41906 128556
rect 41986 128532 41987 128556
rect 42459 128532 42460 128556
rect 42540 128532 42541 128556
rect 43013 128532 43014 128556
rect 43094 128532 43095 128556
rect 43567 128532 43568 128556
rect 43648 128532 43649 128556
rect 44121 128532 44122 128556
rect 44202 128532 44203 128556
rect 44675 128532 44676 128556
rect 44756 128532 44757 128556
rect 45229 128532 45230 128556
rect 45310 128532 45311 128556
rect 45783 128532 45784 128556
rect 45864 128532 45865 128556
rect 46337 128532 46338 128556
rect 46418 128532 46419 128556
rect 46891 128532 46892 128556
rect 46972 128532 46973 128556
rect 47445 128532 47446 128556
rect 47526 128532 47527 128556
rect 47999 128532 48000 128556
rect 48080 128532 48081 128556
rect 48553 128532 48554 128556
rect 48634 128532 48635 128556
rect 49107 128532 49108 128556
rect 49188 128532 49189 128556
rect 49661 128532 49662 128556
rect 49742 128532 49743 128556
rect 50215 128532 50216 128556
rect 50296 128532 50297 128556
rect 50769 128532 50770 128556
rect 50850 128532 50851 128556
rect 51323 128532 51324 128556
rect 51404 128532 51405 128556
rect 40821 128508 40855 128520
rect 41375 128508 41409 128520
rect 41929 128508 41963 128520
rect 42483 128508 42517 128520
rect 43037 128508 43071 128520
rect 43591 128508 43625 128520
rect 44145 128508 44179 128520
rect 44699 128508 44733 128520
rect 45253 128508 45287 128520
rect 45807 128508 45841 128520
rect 46361 128508 46395 128520
rect 46915 128508 46949 128520
rect 47469 128508 47503 128520
rect 48023 128508 48057 128520
rect 48577 128508 48611 128520
rect 49131 128508 49165 128520
rect 49685 128508 49719 128520
rect 50239 128508 50273 128520
rect 50793 128508 50827 128520
rect 51347 128508 51381 128520
rect 2377 127308 2378 127332
rect 2458 127308 2459 127332
rect 2931 127308 2932 127332
rect 3012 127308 3013 127332
rect 3485 127308 3486 127332
rect 3566 127308 3567 127332
rect 4039 127308 4040 127332
rect 4120 127308 4121 127332
rect 4593 127308 4594 127332
rect 4674 127308 4675 127332
rect 5147 127308 5148 127332
rect 5228 127308 5229 127332
rect 5701 127308 5702 127332
rect 5782 127308 5783 127332
rect 6255 127308 6256 127332
rect 6336 127308 6337 127332
rect 6809 127308 6810 127332
rect 6890 127308 6891 127332
rect 7363 127308 7364 127332
rect 7444 127308 7445 127332
rect 7917 127308 7918 127332
rect 7998 127308 7999 127332
rect 8471 127308 8472 127332
rect 8552 127308 8553 127332
rect 9025 127308 9026 127332
rect 9106 127308 9107 127332
rect 9579 127308 9580 127332
rect 9660 127308 9661 127332
rect 10133 127308 10134 127332
rect 10214 127308 10215 127332
rect 10687 127308 10688 127332
rect 10768 127308 10769 127332
rect 11241 127308 11242 127332
rect 11322 127308 11323 127332
rect 11795 127308 11796 127332
rect 11876 127308 11877 127332
rect 12349 127308 12350 127332
rect 12430 127308 12431 127332
rect 2401 127284 2435 127296
rect 2955 127284 2989 127296
rect 3509 127284 3543 127296
rect 4063 127284 4097 127296
rect 4617 127284 4651 127296
rect 5171 127284 5205 127296
rect 5725 127284 5759 127296
rect 6279 127284 6313 127296
rect 6833 127284 6867 127296
rect 7387 127284 7421 127296
rect 7941 127284 7975 127296
rect 8495 127284 8529 127296
rect 9049 127284 9083 127296
rect 9603 127284 9637 127296
rect 10157 127284 10191 127296
rect 10711 127284 10745 127296
rect 11265 127284 11299 127296
rect 11819 127284 11853 127296
rect 12373 127284 12407 127296
rect 2317 125308 2318 125332
rect 2398 125308 2399 125332
rect 3153 125308 3154 125332
rect 3234 125308 3235 125332
rect 3989 125308 3990 125332
rect 4070 125308 4071 125332
rect 4825 125308 4826 125332
rect 4906 125308 4907 125332
rect 5661 125308 5662 125332
rect 5742 125308 5743 125332
rect 6497 125308 6498 125332
rect 6578 125308 6579 125332
rect 7333 125308 7334 125332
rect 7414 125308 7415 125332
rect 8169 125308 8170 125332
rect 8250 125308 8251 125332
rect 9005 125308 9006 125332
rect 9086 125308 9087 125332
rect 9841 125308 9842 125332
rect 9922 125308 9923 125332
rect 10677 125308 10678 125332
rect 10758 125308 10759 125332
rect 11513 125308 11514 125332
rect 11594 125308 11595 125332
rect 12349 125308 12350 125332
rect 12430 125308 12431 125332
rect 2341 125284 2375 125296
rect 3177 125284 3211 125296
rect 4013 125284 4047 125296
rect 4849 125284 4883 125296
rect 5685 125284 5719 125296
rect 6521 125284 6555 125296
rect 7357 125284 7391 125296
rect 8193 125284 8227 125296
rect 9029 125284 9063 125296
rect 9865 125284 9899 125296
rect 10701 125284 10735 125296
rect 11537 125284 11571 125296
rect 12373 125284 12407 125296
rect 22784 124500 22856 128500
rect 23055 124533 23173 128467
rect 23444 124500 23504 128500
rect 23704 124500 23776 128500
rect 23975 124533 24093 128467
rect 24364 124500 24424 128500
rect 24624 124500 24696 128500
rect 24895 124533 25013 128467
rect 25284 124500 25344 128500
rect 25544 124500 25616 128500
rect 25815 124533 25933 128467
rect 26204 124500 26264 128500
rect 26464 124500 26536 128500
rect 26735 124533 26853 128467
rect 27124 124500 27184 128500
rect 27384 124500 27456 128500
rect 27655 124533 27773 128467
rect 28044 124500 28104 128500
rect 28304 124500 28376 128500
rect 28575 124533 28693 128467
rect 28964 124500 29024 128500
rect 29224 124500 29296 128500
rect 29495 124533 29613 128467
rect 29884 124500 29944 128500
rect 30144 124500 30216 128500
rect 30415 124533 30533 128467
rect 30804 124500 30864 128500
rect 31064 124500 31136 128500
rect 31335 124533 31453 128467
rect 31724 124500 31784 128500
rect 31984 124500 32056 128500
rect 32255 124533 32373 128467
rect 32644 124500 32704 128500
rect 59624 127964 59696 129964
rect 59895 127997 60013 129891
rect 60284 127964 60344 129964
rect 60544 127964 60616 129964
rect 60815 127997 60933 129891
rect 61204 127964 61264 129964
rect 61464 127964 61536 129964
rect 61735 127997 61853 129891
rect 62124 127964 62184 129964
rect 62384 127964 62456 129964
rect 62655 127997 62773 129891
rect 63044 127964 63104 129964
rect 63304 127964 63376 129964
rect 63575 127997 63693 129891
rect 63964 127964 64024 129964
rect 64224 127964 64296 129964
rect 64495 127997 64613 129891
rect 64884 127964 64944 129964
rect 65144 127964 65216 129964
rect 65415 127997 65533 129891
rect 65804 127964 65864 129964
rect 66064 127964 66136 129964
rect 66335 127997 66453 129891
rect 66724 127964 66784 129964
rect 66984 127964 67056 129964
rect 67255 127997 67373 129891
rect 67644 127964 67704 129964
rect 67904 127964 67976 129964
rect 68175 127997 68293 129891
rect 68564 127964 68624 129964
rect 68824 127964 68896 129964
rect 69095 127997 69213 129891
rect 69484 127964 69544 129964
rect 80176 128934 80248 130934
rect 80447 128967 80565 130861
rect 80836 128934 80896 130934
rect 81096 128934 81168 130934
rect 81367 128967 81485 130861
rect 81756 128934 81816 130934
rect 82016 128934 82088 130934
rect 82287 128967 82405 130861
rect 82676 128934 82736 130934
rect 82936 128934 83008 130934
rect 83207 128967 83325 130861
rect 83596 128934 83656 130934
rect 83856 128934 83928 130934
rect 84127 128967 84245 130861
rect 84516 128934 84576 130934
rect 84776 128934 84848 130934
rect 85047 128967 85165 130861
rect 85436 128934 85496 130934
rect 85696 128934 85768 130934
rect 85967 128967 86085 130861
rect 86356 128934 86416 130934
rect 86616 128934 86688 130934
rect 86887 128967 87005 130861
rect 87276 128934 87336 130934
rect 87536 128934 87608 130934
rect 87807 128967 87925 130861
rect 88196 128934 88256 130934
rect 88456 128934 88528 130934
rect 88727 128967 88845 130861
rect 89116 128934 89176 130934
rect 89376 128934 89448 130934
rect 89647 128967 89765 130861
rect 90036 128934 90096 130934
rect 121650 130927 121653 130928
rect 121650 130926 121651 130927
rect 121652 130926 121653 130927
rect 121650 130925 121653 130926
rect 119603 130817 121521 130899
rect 133592 130823 134592 130951
rect 121650 130790 121653 130791
rect 121650 130789 121651 130790
rect 121652 130789 121653 130790
rect 121650 130788 121653 130789
rect 99739 129696 99740 129720
rect 99820 129696 99821 129720
rect 100293 129696 100294 129720
rect 100374 129696 100375 129720
rect 100847 129696 100848 129720
rect 100928 129696 100929 129720
rect 101401 129696 101402 129720
rect 101482 129696 101483 129720
rect 101955 129696 101956 129720
rect 102036 129696 102037 129720
rect 102509 129696 102510 129720
rect 102590 129696 102591 129720
rect 103063 129696 103064 129720
rect 103144 129696 103145 129720
rect 103617 129696 103618 129720
rect 103698 129696 103699 129720
rect 104171 129696 104172 129720
rect 104252 129696 104253 129720
rect 104725 129696 104726 129720
rect 104806 129696 104807 129720
rect 105279 129696 105280 129720
rect 105360 129696 105361 129720
rect 105833 129696 105834 129720
rect 105914 129696 105915 129720
rect 106387 129696 106388 129720
rect 106468 129696 106469 129720
rect 106941 129696 106942 129720
rect 107022 129696 107023 129720
rect 107495 129696 107496 129720
rect 107576 129696 107577 129720
rect 108049 129696 108050 129720
rect 108130 129696 108131 129720
rect 108603 129696 108604 129720
rect 108684 129696 108685 129720
rect 109157 129696 109158 129720
rect 109238 129696 109239 129720
rect 109711 129696 109712 129720
rect 109792 129696 109793 129720
rect 110265 129696 110266 129720
rect 110346 129696 110347 129720
rect 99763 129672 99797 129684
rect 100317 129672 100351 129684
rect 100871 129672 100905 129684
rect 101425 129672 101459 129684
rect 101979 129672 102013 129684
rect 102533 129672 102567 129684
rect 103087 129672 103121 129684
rect 103641 129672 103675 129684
rect 104195 129672 104229 129684
rect 104749 129672 104783 129684
rect 105303 129672 105337 129684
rect 105857 129672 105891 129684
rect 106411 129672 106445 129684
rect 106965 129672 106999 129684
rect 107519 129672 107553 129684
rect 108073 129672 108107 129684
rect 108627 129672 108661 129684
rect 109181 129672 109215 129684
rect 109735 129672 109769 129684
rect 110289 129672 110323 129684
rect 119390 129681 119472 130715
rect 119682 129851 119764 130545
rect 119904 130532 121210 130614
rect 120072 130350 121014 130400
rect 119941 130299 119967 130310
rect 119957 130259 120051 130299
rect 120963 130259 121057 130299
rect 119957 130099 120051 130139
rect 120963 130099 121057 130139
rect 119941 130088 119967 130099
rect 120072 130006 121014 130056
rect 119904 129780 121210 129862
rect 121250 129851 121332 130545
rect 121542 129681 121624 130715
rect 127486 130689 128486 130739
rect 128882 130689 129482 130739
rect 127486 130533 128486 130661
rect 131226 130629 132226 130679
rect 133592 130673 134592 130723
rect 128882 130533 129482 130589
rect 127486 130377 128486 130505
rect 128882 130377 129482 130433
rect 131226 130413 132226 130541
rect 127486 130227 128486 130277
rect 128882 130221 129482 130277
rect 131226 130203 132226 130253
rect 128882 130071 129482 130121
rect 119603 129498 121521 129580
rect 120316 129443 120486 129498
rect 121550 129443 121719 129511
rect 120384 129363 120385 129443
rect 120418 129403 120486 129443
rect 120418 129363 120485 129403
rect 120384 129362 120485 129363
rect 121618 129363 121619 129443
rect 121652 129363 121719 129443
rect 121618 129362 121719 129363
rect 120693 129142 121293 129192
rect 120693 128892 121293 128942
rect 122413 128467 122463 129467
rect 122623 128467 122751 129467
rect 122839 128467 122967 129467
rect 123055 128467 123183 129467
rect 123271 128467 123399 129467
rect 123487 128467 123543 129467
rect 123703 128467 123759 129467
rect 123919 128467 124047 129467
rect 124135 128467 124263 129467
rect 124351 128467 124479 129467
rect 124567 128467 124695 129467
rect 124783 128467 124839 129467
rect 124999 128467 125127 129467
rect 125215 128467 125343 129467
rect 125431 128467 125559 129467
rect 125647 128467 125697 129467
rect 125763 128467 125813 129467
rect 125973 128467 126023 129467
rect 126089 128467 126139 129467
rect 126299 128467 126349 129467
rect 126415 128467 126465 129467
rect 126625 128467 126675 129467
rect 126738 129282 126750 129482
rect 126741 128467 126791 129067
rect 126991 128467 127047 129067
rect 127147 128467 127275 129067
rect 127303 128467 127359 129067
rect 127459 128467 127587 129067
rect 127615 128467 127665 129067
rect 127731 128467 127781 129467
rect 127881 128467 127937 129467
rect 128037 128467 128087 129467
rect 128165 128467 128215 129467
rect 128315 128467 128443 129467
rect 128471 128467 128599 129467
rect 128627 128467 128683 129467
rect 128783 128467 128911 129467
rect 128939 128467 129067 129467
rect 129095 128467 129223 129467
rect 129251 128467 129301 129467
rect 129367 128467 129417 129467
rect 129517 128467 129645 129467
rect 129673 128467 129801 129467
rect 129829 128467 129957 129467
rect 129985 128467 130041 129467
rect 130141 128467 130269 129467
rect 130297 128467 130425 129467
rect 130453 128467 130509 129467
rect 130609 128467 130659 129467
rect 131880 129267 131933 129467
rect 131883 128467 131933 129267
rect 132093 128467 132221 129467
rect 132309 128467 132365 129467
rect 132525 128467 132653 129467
rect 132741 128467 132791 129467
rect 132857 128467 132907 129467
rect 133067 128467 133117 129467
rect 130604 128380 130640 128391
rect 130756 128380 133080 128391
rect 130604 128358 133080 128380
rect 130604 128357 130640 128358
rect 130756 128357 133080 128358
rect 41351 126532 41352 126556
rect 41432 126532 41433 126556
rect 41905 126532 41906 126556
rect 41986 126532 41987 126556
rect 42459 126532 42460 126556
rect 42540 126532 42541 126556
rect 43013 126532 43014 126556
rect 43094 126532 43095 126556
rect 43567 126532 43568 126556
rect 43648 126532 43649 126556
rect 44121 126532 44122 126556
rect 44202 126532 44203 126556
rect 44675 126532 44676 126556
rect 44756 126532 44757 126556
rect 45229 126532 45230 126556
rect 45310 126532 45311 126556
rect 45783 126532 45784 126556
rect 45864 126532 45865 126556
rect 46337 126532 46338 126556
rect 46418 126532 46419 126556
rect 46891 126532 46892 126556
rect 46972 126532 46973 126556
rect 47445 126532 47446 126556
rect 47526 126532 47527 126556
rect 47999 126532 48000 126556
rect 48080 126532 48081 126556
rect 48553 126532 48554 126556
rect 48634 126532 48635 126556
rect 49107 126532 49108 126556
rect 49188 126532 49189 126556
rect 49661 126532 49662 126556
rect 49742 126532 49743 126556
rect 50215 126532 50216 126556
rect 50296 126532 50297 126556
rect 50769 126532 50770 126556
rect 50850 126532 50851 126556
rect 51323 126532 51324 126556
rect 51404 126532 51405 126556
rect 41375 126508 41409 126520
rect 41929 126508 41963 126520
rect 42483 126508 42517 126520
rect 43037 126508 43071 126520
rect 43591 126508 43625 126520
rect 44145 126508 44179 126520
rect 44699 126508 44733 126520
rect 45253 126508 45287 126520
rect 45807 126508 45841 126520
rect 46361 126508 46395 126520
rect 46915 126508 46949 126520
rect 47469 126508 47503 126520
rect 48023 126508 48057 126520
rect 48577 126508 48611 126520
rect 49131 126508 49165 126520
rect 49685 126508 49719 126520
rect 50239 126508 50273 126520
rect 50793 126508 50827 126520
rect 51347 126508 51381 126520
rect 41291 124532 41292 124556
rect 41372 124532 41373 124556
rect 42127 124532 42128 124556
rect 42208 124532 42209 124556
rect 42963 124532 42964 124556
rect 43044 124532 43045 124556
rect 43799 124532 43800 124556
rect 43880 124532 43881 124556
rect 44635 124532 44636 124556
rect 44716 124532 44717 124556
rect 45471 124532 45472 124556
rect 45552 124532 45553 124556
rect 46307 124532 46308 124556
rect 46388 124532 46389 124556
rect 47143 124532 47144 124556
rect 47224 124532 47225 124556
rect 47979 124532 47980 124556
rect 48060 124532 48061 124556
rect 48815 124532 48816 124556
rect 48896 124532 48897 124556
rect 49651 124532 49652 124556
rect 49732 124532 49733 124556
rect 50487 124532 50488 124556
rect 50568 124532 50569 124556
rect 51323 124532 51324 124556
rect 51404 124532 51405 124556
rect 41315 124508 41349 124520
rect 42151 124508 42185 124520
rect 42987 124508 43021 124520
rect 43823 124508 43857 124520
rect 44659 124508 44693 124520
rect 45495 124508 45529 124520
rect 46331 124508 46365 124520
rect 47167 124508 47201 124520
rect 48003 124508 48037 124520
rect 48839 124508 48873 124520
rect 49675 124508 49709 124520
rect 50511 124508 50545 124520
rect 51347 124508 51381 124520
rect 2317 123308 2318 123332
rect 2398 123308 2399 123332
rect 3153 123308 3154 123332
rect 3234 123308 3235 123332
rect 3989 123308 3990 123332
rect 4070 123308 4071 123332
rect 4825 123308 4826 123332
rect 4906 123308 4907 123332
rect 5661 123308 5662 123332
rect 5742 123308 5743 123332
rect 6497 123308 6498 123332
rect 6578 123308 6579 123332
rect 7333 123308 7334 123332
rect 7414 123308 7415 123332
rect 8169 123308 8170 123332
rect 8250 123308 8251 123332
rect 9005 123308 9006 123332
rect 9086 123308 9087 123332
rect 9841 123308 9842 123332
rect 9922 123308 9923 123332
rect 10677 123308 10678 123332
rect 10758 123308 10759 123332
rect 11513 123308 11514 123332
rect 11594 123308 11595 123332
rect 12349 123308 12350 123332
rect 12430 123308 12431 123332
rect 2341 123284 2375 123296
rect 3177 123284 3211 123296
rect 4013 123284 4047 123296
rect 4849 123284 4883 123296
rect 5685 123284 5719 123296
rect 6521 123284 6555 123296
rect 7357 123284 7391 123296
rect 8193 123284 8227 123296
rect 9029 123284 9063 123296
rect 9865 123284 9899 123296
rect 10701 123284 10735 123296
rect 11537 123284 11571 123296
rect 12373 123284 12407 123296
rect 2317 121308 2318 121332
rect 2398 121308 2399 121332
rect 3153 121308 3154 121332
rect 3234 121308 3235 121332
rect 3989 121308 3990 121332
rect 4070 121308 4071 121332
rect 4825 121308 4826 121332
rect 4906 121308 4907 121332
rect 5661 121308 5662 121332
rect 5742 121308 5743 121332
rect 6497 121308 6498 121332
rect 6578 121308 6579 121332
rect 7333 121308 7334 121332
rect 7414 121308 7415 121332
rect 8169 121308 8170 121332
rect 8250 121308 8251 121332
rect 9005 121308 9006 121332
rect 9086 121308 9087 121332
rect 9841 121308 9842 121332
rect 9922 121308 9923 121332
rect 10677 121308 10678 121332
rect 10758 121308 10759 121332
rect 11513 121308 11514 121332
rect 11594 121308 11595 121332
rect 12349 121308 12350 121332
rect 12430 121308 12431 121332
rect 2341 121284 2375 121296
rect 3177 121284 3211 121296
rect 4013 121284 4047 121296
rect 4849 121284 4883 121296
rect 5685 121284 5719 121296
rect 6521 121284 6555 121296
rect 7357 121284 7391 121296
rect 8193 121284 8227 121296
rect 9029 121284 9063 121296
rect 9865 121284 9899 121296
rect 10701 121284 10735 121296
rect 11537 121284 11571 121296
rect 12373 121284 12407 121296
rect 22784 119900 22856 123900
rect 23055 119933 23173 123867
rect 23444 119900 23504 123900
rect 23704 119900 23776 123900
rect 23975 119933 24093 123867
rect 24364 119900 24424 123900
rect 24624 119900 24696 123900
rect 24895 119933 25013 123867
rect 25284 119900 25344 123900
rect 25544 119900 25616 123900
rect 25815 119933 25933 123867
rect 26204 119900 26264 123900
rect 26464 119900 26536 123900
rect 26735 119933 26853 123867
rect 27124 119900 27184 123900
rect 27384 119900 27456 123900
rect 27655 119933 27773 123867
rect 28044 119900 28104 123900
rect 28304 119900 28376 123900
rect 28575 119933 28693 123867
rect 28964 119900 29024 123900
rect 29224 119900 29296 123900
rect 29495 119933 29613 123867
rect 29884 119900 29944 123900
rect 30144 119900 30216 123900
rect 30415 119933 30533 123867
rect 30804 119900 30864 123900
rect 31064 119900 31136 123900
rect 31335 119933 31453 123867
rect 31724 119900 31784 123900
rect 31984 119900 32056 123900
rect 32255 119933 32373 123867
rect 32644 119900 32704 123900
rect 59624 123364 59696 127364
rect 59895 123397 60013 127331
rect 60284 123364 60344 127364
rect 60544 123364 60616 127364
rect 60815 123397 60933 127331
rect 61204 123364 61264 127364
rect 61464 123364 61536 127364
rect 61735 123397 61853 127331
rect 62124 123364 62184 127364
rect 62384 123364 62456 127364
rect 62655 123397 62773 127331
rect 63044 123364 63104 127364
rect 63304 123364 63376 127364
rect 63575 123397 63693 127331
rect 63964 123364 64024 127364
rect 64224 123364 64296 127364
rect 64495 123397 64613 127331
rect 64884 123364 64944 127364
rect 65144 123364 65216 127364
rect 65415 123397 65533 127331
rect 65804 123364 65864 127364
rect 66064 123364 66136 127364
rect 66335 123397 66453 127331
rect 66724 123364 66784 127364
rect 66984 123364 67056 127364
rect 67255 123397 67373 127331
rect 67644 123364 67704 127364
rect 67904 123364 67976 127364
rect 68175 123397 68293 127331
rect 68564 123364 68624 127364
rect 68824 123364 68896 127364
rect 69095 123397 69213 127331
rect 69484 123364 69544 127364
rect 80176 124334 80248 128334
rect 80447 124367 80565 128301
rect 80836 124334 80896 128334
rect 81096 124334 81168 128334
rect 81367 124367 81485 128301
rect 81756 124334 81816 128334
rect 82016 124334 82088 128334
rect 82287 124367 82405 128301
rect 82676 124334 82736 128334
rect 82936 124334 83008 128334
rect 83207 124367 83325 128301
rect 83596 124334 83656 128334
rect 83856 124334 83928 128334
rect 84127 124367 84245 128301
rect 84516 124334 84576 128334
rect 84776 124334 84848 128334
rect 85047 124367 85165 128301
rect 85436 124334 85496 128334
rect 85696 124334 85768 128334
rect 85967 124367 86085 128301
rect 86356 124334 86416 128334
rect 86616 124334 86688 128334
rect 86887 124367 87005 128301
rect 87276 124334 87336 128334
rect 87536 124334 87608 128334
rect 87807 124367 87925 128301
rect 88196 124334 88256 128334
rect 88456 124334 88528 128334
rect 88727 124367 88845 128301
rect 89116 124334 89176 128334
rect 89376 124334 89448 128334
rect 89647 124367 89765 128301
rect 90036 124334 90096 128334
rect 100293 127696 100294 127720
rect 100374 127696 100375 127720
rect 100847 127696 100848 127720
rect 100928 127696 100929 127720
rect 101401 127696 101402 127720
rect 101482 127696 101483 127720
rect 101955 127696 101956 127720
rect 102036 127696 102037 127720
rect 102509 127696 102510 127720
rect 102590 127696 102591 127720
rect 103063 127696 103064 127720
rect 103144 127696 103145 127720
rect 103617 127696 103618 127720
rect 103698 127696 103699 127720
rect 104171 127696 104172 127720
rect 104252 127696 104253 127720
rect 104725 127696 104726 127720
rect 104806 127696 104807 127720
rect 105279 127696 105280 127720
rect 105360 127696 105361 127720
rect 105833 127696 105834 127720
rect 105914 127696 105915 127720
rect 106387 127696 106388 127720
rect 106468 127696 106469 127720
rect 106941 127696 106942 127720
rect 107022 127696 107023 127720
rect 107495 127696 107496 127720
rect 107576 127696 107577 127720
rect 108049 127696 108050 127720
rect 108130 127696 108131 127720
rect 108603 127696 108604 127720
rect 108684 127696 108685 127720
rect 109157 127696 109158 127720
rect 109238 127696 109239 127720
rect 109711 127696 109712 127720
rect 109792 127696 109793 127720
rect 110265 127696 110266 127720
rect 110346 127696 110347 127720
rect 100317 127672 100351 127684
rect 100871 127672 100905 127684
rect 101425 127672 101459 127684
rect 101979 127672 102013 127684
rect 102533 127672 102567 127684
rect 103087 127672 103121 127684
rect 103641 127672 103675 127684
rect 104195 127672 104229 127684
rect 104749 127672 104783 127684
rect 105303 127672 105337 127684
rect 105857 127672 105891 127684
rect 106411 127672 106445 127684
rect 106965 127672 106999 127684
rect 107519 127672 107553 127684
rect 108073 127672 108107 127684
rect 108627 127672 108661 127684
rect 109181 127672 109215 127684
rect 109735 127672 109769 127684
rect 110289 127672 110323 127684
rect 125666 127148 125736 127180
rect 125770 127148 125805 127180
rect 125839 127148 125874 127180
rect 125908 127148 125942 127180
rect 125976 127148 126010 127180
rect 126044 127148 126078 127180
rect 126112 127148 126146 127180
rect 126180 127148 126214 127180
rect 126248 127148 126282 127180
rect 126316 127148 126350 127180
rect 126384 127148 126418 127180
rect 126452 127148 126486 127180
rect 126520 127148 126554 127180
rect 126588 127148 126622 127180
rect 126656 127148 126690 127180
rect 126724 127148 126758 127180
rect 126792 127148 126826 127180
rect 126860 127148 126894 127180
rect 126928 127148 126962 127180
rect 126996 127148 127030 127180
rect 127064 127148 127098 127180
rect 127132 127148 127166 127180
rect 127200 127148 127234 127180
rect 127268 127148 127302 127180
rect 127336 127148 127370 127180
rect 127404 127148 127438 127180
rect 127472 127148 127506 127180
rect 127540 127148 127574 127180
rect 127608 127148 127642 127180
rect 127676 127148 127710 127180
rect 127744 127148 127778 127180
rect 127812 127148 127846 127180
rect 127880 127148 127914 127180
rect 127948 127148 127982 127180
rect 128016 127148 128050 127180
rect 128084 127148 128118 127180
rect 128152 127148 128186 127180
rect 128220 127148 128254 127180
rect 128288 127148 128322 127180
rect 128356 127148 128390 127180
rect 128424 127148 128458 127180
rect 128492 127148 128526 127180
rect 128560 127148 128594 127180
rect 128628 127148 128662 127180
rect 128696 127148 128730 127180
rect 128764 127148 128798 127180
rect 128832 127148 128866 127180
rect 128900 127148 128934 127180
rect 128968 127148 129002 127180
rect 129036 127148 129070 127180
rect 129104 127148 129138 127180
rect 129172 127148 129206 127180
rect 129240 127148 129274 127180
rect 129308 127148 129342 127180
rect 129376 127148 129410 127180
rect 129444 127148 129478 127180
rect 129512 127148 129546 127180
rect 129580 127148 129614 127180
rect 129648 127148 129682 127180
rect 129716 127148 129750 127180
rect 129784 127148 129818 127180
rect 129852 127148 129886 127180
rect 129920 127148 129954 127180
rect 129988 127148 130022 127180
rect 130056 127148 130090 127180
rect 130124 127148 130158 127180
rect 130192 127148 130226 127180
rect 130260 127148 130294 127180
rect 130328 127148 130362 127180
rect 130396 127148 130430 127180
rect 130464 127148 130498 127180
rect 130532 127148 130566 127180
rect 130600 127148 130634 127180
rect 130668 127148 130702 127180
rect 130736 127148 130770 127180
rect 130804 127148 130838 127180
rect 130872 127148 130906 127180
rect 130940 127148 130974 127180
rect 131008 127148 131042 127180
rect 131076 127148 131110 127180
rect 131144 127148 131178 127180
rect 131212 127148 131246 127180
rect 131280 127148 131314 127180
rect 131348 127148 131382 127180
rect 131416 127148 131450 127180
rect 131484 127148 131518 127180
rect 131552 127148 131586 127180
rect 131620 127148 131654 127180
rect 131688 127148 131722 127180
rect 131756 127148 131790 127180
rect 131824 127148 131858 127180
rect 131892 127148 131926 127180
rect 131960 127148 131994 127180
rect 132028 127148 132062 127180
rect 132096 127148 132130 127180
rect 132164 127148 132198 127180
rect 132232 127148 132266 127180
rect 132300 127148 132334 127180
rect 132368 127148 132402 127180
rect 132436 127148 132470 127180
rect 132504 127148 132538 127180
rect 132572 127148 132606 127180
rect 132640 127148 132680 127180
rect 132777 127148 132848 127216
rect 134612 127174 134626 127180
rect 125736 127126 125770 127148
rect 125805 127126 125839 127148
rect 125874 127126 125908 127148
rect 125942 127126 125976 127148
rect 126010 127126 126044 127148
rect 126078 127126 126112 127148
rect 126146 127126 126180 127148
rect 126214 127126 126248 127148
rect 126282 127126 126316 127148
rect 126350 127126 126384 127148
rect 126418 127126 126452 127148
rect 126486 127126 126520 127148
rect 126554 127126 126588 127148
rect 126622 127126 126656 127148
rect 126690 127126 126724 127148
rect 126758 127126 126792 127148
rect 126826 127126 126860 127148
rect 126894 127126 126928 127148
rect 126962 127126 126996 127148
rect 127030 127126 127064 127148
rect 127098 127126 127132 127148
rect 127166 127126 127200 127148
rect 127234 127126 127268 127148
rect 127302 127126 127336 127148
rect 127370 127126 127404 127148
rect 127438 127126 127472 127148
rect 127506 127126 127540 127148
rect 127574 127126 127608 127148
rect 127642 127126 127676 127148
rect 127710 127126 127744 127148
rect 127778 127126 127812 127148
rect 127846 127126 127880 127148
rect 127914 127126 127948 127148
rect 127982 127126 128016 127148
rect 128050 127126 128084 127148
rect 128118 127126 128152 127148
rect 128186 127126 128220 127148
rect 128254 127126 128288 127148
rect 128322 127126 128356 127148
rect 128390 127126 128424 127148
rect 128458 127126 128492 127148
rect 128526 127126 128560 127148
rect 128594 127126 128628 127148
rect 128662 127126 128696 127148
rect 128730 127126 128764 127148
rect 128798 127126 128832 127148
rect 128866 127126 128900 127148
rect 128934 127126 128968 127148
rect 129002 127126 129036 127148
rect 129070 127126 129104 127148
rect 129138 127126 129172 127148
rect 129206 127126 129240 127148
rect 129274 127126 129308 127148
rect 129342 127126 129376 127148
rect 129410 127126 129444 127148
rect 129478 127126 129512 127148
rect 129546 127126 129580 127148
rect 129614 127126 129648 127148
rect 129682 127126 129716 127148
rect 129750 127126 129784 127148
rect 129818 127126 129852 127148
rect 129886 127126 129920 127148
rect 129954 127126 129988 127148
rect 130022 127126 130056 127148
rect 130090 127126 130124 127148
rect 130158 127126 130192 127148
rect 130226 127126 130260 127148
rect 130294 127126 130328 127148
rect 130362 127126 130396 127148
rect 130430 127126 130464 127148
rect 130498 127126 130532 127148
rect 130566 127126 130600 127148
rect 130634 127126 130668 127148
rect 130702 127126 130736 127148
rect 130770 127126 130804 127148
rect 130838 127126 130872 127148
rect 130906 127126 130940 127148
rect 130974 127126 131008 127148
rect 131042 127126 131076 127148
rect 131110 127126 131144 127148
rect 131178 127126 131212 127148
rect 131246 127126 131280 127148
rect 131314 127126 131348 127148
rect 131382 127126 131416 127148
rect 131450 127126 131484 127148
rect 131518 127126 131552 127148
rect 131586 127126 131620 127148
rect 131654 127126 131688 127148
rect 131722 127126 131756 127148
rect 131790 127126 131824 127148
rect 131858 127126 131892 127148
rect 131926 127126 131960 127148
rect 131994 127126 132028 127148
rect 132062 127126 132096 127148
rect 132130 127126 132164 127148
rect 132198 127126 132232 127148
rect 132266 127126 132300 127148
rect 132334 127126 132368 127148
rect 132402 127126 132436 127148
rect 132470 127126 132504 127148
rect 132538 127126 132572 127148
rect 132606 127126 132640 127148
rect 132680 127127 132777 127148
rect 132780 127127 132848 127148
rect 132680 127126 132848 127127
rect 125666 127094 132680 127126
rect 120992 126779 121992 126829
rect 122102 126779 123102 126829
rect 123223 126779 124223 126829
rect 124344 126779 125344 126829
rect 125901 126779 126901 126829
rect 127022 126779 128022 126829
rect 128143 126779 129143 126829
rect 129253 126779 130253 126829
rect 130374 126779 131374 126829
rect 131495 126779 132495 126829
rect 120992 126609 121992 126659
rect 122102 126609 123102 126659
rect 123223 126609 124223 126659
rect 124344 126609 125344 126659
rect 125901 126609 126901 126659
rect 127022 126609 128022 126659
rect 128143 126609 129143 126659
rect 129253 126609 130253 126659
rect 130374 126609 131374 126659
rect 131495 126609 132495 126659
rect 132777 126350 132848 126380
rect 134572 126350 134612 127174
rect 120597 126346 120732 126350
rect 125606 126346 125640 126350
rect 120597 126312 132680 126346
rect 132777 126336 134612 126350
rect 132777 126322 134602 126336
rect 132777 126312 132848 126322
rect 120596 126296 120597 126312
rect 132680 126297 132777 126312
rect 132780 126297 132848 126312
rect 132680 126296 132848 126297
rect 134626 126296 134666 127174
rect 120597 126258 132680 126296
rect 132820 126282 134666 126296
rect 132820 126268 134656 126282
rect 100233 125696 100234 125720
rect 100314 125696 100315 125720
rect 101069 125696 101070 125720
rect 101150 125696 101151 125720
rect 101905 125696 101906 125720
rect 101986 125696 101987 125720
rect 102741 125696 102742 125720
rect 102822 125696 102823 125720
rect 103577 125696 103578 125720
rect 103658 125696 103659 125720
rect 104413 125696 104414 125720
rect 104494 125696 104495 125720
rect 105249 125696 105250 125720
rect 105330 125696 105331 125720
rect 106085 125696 106086 125720
rect 106166 125696 106167 125720
rect 106921 125696 106922 125720
rect 107002 125696 107003 125720
rect 107757 125696 107758 125720
rect 107838 125696 107839 125720
rect 108593 125696 108594 125720
rect 108674 125696 108675 125720
rect 109429 125696 109430 125720
rect 109510 125696 109511 125720
rect 110265 125696 110266 125720
rect 110346 125696 110347 125720
rect 100257 125672 100291 125684
rect 101093 125672 101127 125684
rect 101929 125672 101963 125684
rect 102765 125672 102799 125684
rect 103601 125672 103635 125684
rect 104437 125672 104471 125684
rect 105273 125672 105307 125684
rect 106109 125672 106143 125684
rect 106945 125672 106979 125684
rect 107781 125672 107815 125684
rect 108617 125672 108651 125684
rect 109453 125672 109487 125684
rect 110289 125672 110323 125684
rect 121219 124928 121429 124964
rect 133481 124928 133594 124964
rect 134043 124928 134325 124964
rect 120808 123928 120886 124928
rect 121008 123928 121080 124928
rect 121231 123928 121255 124928
rect 121296 123928 121352 124928
rect 121393 123928 121429 124928
rect 121654 123928 121714 124928
rect 121914 123928 121986 124928
rect 122216 123928 122272 124928
rect 122288 123928 122344 124928
rect 122646 123928 122706 124928
rect 122906 123928 122978 124928
rect 123208 123928 123264 124928
rect 123280 123928 123336 124928
rect 123638 123928 123698 124928
rect 123898 123928 123970 124928
rect 124200 123928 124256 124928
rect 124272 123928 124328 124928
rect 124630 123928 124690 124928
rect 124890 123928 124962 124928
rect 125192 123928 125248 124928
rect 125264 123928 125320 124928
rect 125622 123928 125682 124928
rect 125882 123928 125954 124928
rect 126184 123928 126240 124928
rect 126256 123928 126312 124928
rect 126614 123928 126674 124928
rect 126874 123928 126946 124928
rect 127176 123928 127232 124928
rect 127248 123928 127304 124928
rect 127606 123928 127666 124928
rect 127866 123928 127938 124928
rect 128168 123928 128224 124928
rect 128240 123928 128296 124928
rect 128598 123928 128658 124928
rect 128858 123928 128930 124928
rect 129160 123928 129216 124928
rect 129232 123928 129288 124928
rect 129590 123928 129650 124928
rect 129850 123928 129922 124928
rect 130152 123928 130208 124928
rect 130224 123928 130280 124928
rect 130582 123928 130642 124928
rect 130842 123928 130914 124928
rect 131144 123928 131200 124928
rect 131216 123928 131272 124928
rect 131574 123928 131634 124928
rect 131834 123928 131906 124928
rect 132136 123928 132192 124928
rect 132208 123928 132264 124928
rect 132566 123928 132626 124928
rect 132826 123928 132898 124928
rect 133128 123928 133184 124928
rect 133200 123928 133256 124928
rect 133481 123928 133517 124928
rect 133558 123928 133594 124928
rect 133818 123928 133890 124928
rect 134043 123928 134079 124928
rect 134120 123928 134176 124928
rect 134192 123928 134248 124928
rect 134289 123928 134325 124928
rect 134536 123928 134596 124928
rect 134632 123928 134736 124928
rect 140710 124063 140788 125063
rect 140910 124063 140982 125063
rect 161216 124211 161280 124247
rect 121219 123892 121429 123928
rect 133481 123892 133594 123928
rect 134043 123892 134325 123928
rect 41291 122532 41292 122556
rect 41372 122532 41373 122556
rect 42127 122532 42128 122556
rect 42208 122532 42209 122556
rect 42963 122532 42964 122556
rect 43044 122532 43045 122556
rect 43799 122532 43800 122556
rect 43880 122532 43881 122556
rect 44635 122532 44636 122556
rect 44716 122532 44717 122556
rect 45471 122532 45472 122556
rect 45552 122532 45553 122556
rect 46307 122532 46308 122556
rect 46388 122532 46389 122556
rect 47143 122532 47144 122556
rect 47224 122532 47225 122556
rect 47979 122532 47980 122556
rect 48060 122532 48061 122556
rect 48815 122532 48816 122556
rect 48896 122532 48897 122556
rect 49651 122532 49652 122556
rect 49732 122532 49733 122556
rect 50487 122532 50488 122556
rect 50568 122532 50569 122556
rect 51323 122532 51324 122556
rect 51404 122532 51405 122556
rect 41315 122508 41349 122520
rect 42151 122508 42185 122520
rect 42987 122508 43021 122520
rect 43823 122508 43857 122520
rect 44659 122508 44693 122520
rect 45495 122508 45529 122520
rect 46331 122508 46365 122520
rect 47167 122508 47201 122520
rect 48003 122508 48037 122520
rect 48839 122508 48873 122520
rect 49675 122508 49709 122520
rect 50511 122508 50545 122520
rect 51347 122508 51381 122520
rect 41291 120532 41292 120556
rect 41372 120532 41373 120556
rect 42127 120532 42128 120556
rect 42208 120532 42209 120556
rect 42963 120532 42964 120556
rect 43044 120532 43045 120556
rect 43799 120532 43800 120556
rect 43880 120532 43881 120556
rect 44635 120532 44636 120556
rect 44716 120532 44717 120556
rect 45471 120532 45472 120556
rect 45552 120532 45553 120556
rect 46307 120532 46308 120556
rect 46388 120532 46389 120556
rect 47143 120532 47144 120556
rect 47224 120532 47225 120556
rect 47979 120532 47980 120556
rect 48060 120532 48061 120556
rect 48815 120532 48816 120556
rect 48896 120532 48897 120556
rect 49651 120532 49652 120556
rect 49732 120532 49733 120556
rect 50487 120532 50488 120556
rect 50568 120532 50569 120556
rect 51323 120532 51324 120556
rect 51404 120532 51405 120556
rect 41315 120508 41349 120520
rect 42151 120508 42185 120520
rect 42987 120508 43021 120520
rect 43823 120508 43857 120520
rect 44659 120508 44693 120520
rect 45495 120508 45529 120520
rect 46331 120508 46365 120520
rect 47167 120508 47201 120520
rect 48003 120508 48037 120520
rect 48839 120508 48873 120520
rect 49675 120508 49709 120520
rect 50511 120508 50545 120520
rect 51347 120508 51381 120520
rect 3989 119308 3990 119332
rect 4070 119308 4071 119332
rect 4825 119308 4826 119332
rect 4906 119308 4907 119332
rect 5661 119308 5662 119332
rect 5742 119308 5743 119332
rect 6497 119308 6498 119332
rect 6578 119308 6579 119332
rect 7333 119308 7334 119332
rect 7414 119308 7415 119332
rect 8169 119308 8170 119332
rect 8250 119308 8251 119332
rect 9005 119308 9006 119332
rect 9086 119308 9087 119332
rect 9841 119308 9842 119332
rect 9922 119308 9923 119332
rect 10677 119308 10678 119332
rect 10758 119308 10759 119332
rect 11513 119308 11514 119332
rect 11594 119308 11595 119332
rect 12349 119308 12350 119332
rect 12430 119308 12431 119332
rect 4013 119284 4047 119296
rect 4849 119284 4883 119296
rect 5685 119284 5719 119296
rect 6521 119284 6555 119296
rect 7357 119284 7391 119296
rect 8193 119284 8227 119296
rect 9029 119284 9063 119296
rect 9865 119284 9899 119296
rect 10701 119284 10735 119296
rect 11537 119284 11571 119296
rect 12373 119284 12407 119296
rect 3989 117687 3990 117711
rect 4070 117687 4071 117711
rect 4825 117687 4826 117711
rect 4906 117687 4907 117711
rect 5661 117687 5662 117711
rect 5742 117687 5743 117711
rect 6497 117687 6498 117711
rect 6578 117687 6579 117711
rect 7333 117687 7334 117711
rect 7414 117687 7415 117711
rect 8169 117687 8170 117711
rect 8250 117687 8251 117711
rect 9005 117687 9006 117711
rect 9086 117687 9087 117711
rect 9841 117687 9842 117711
rect 9922 117687 9923 117711
rect 10677 117687 10678 117711
rect 10758 117687 10759 117711
rect 11513 117687 11514 117711
rect 11594 117687 11595 117711
rect 12349 117687 12350 117711
rect 12430 117687 12431 117711
rect 4013 117663 4047 117675
rect 4849 117663 4883 117675
rect 5685 117663 5719 117675
rect 6521 117663 6555 117675
rect 7357 117663 7391 117675
rect 8193 117663 8227 117675
rect 9029 117663 9063 117675
rect 9865 117663 9899 117675
rect 10701 117663 10735 117675
rect 11537 117663 11571 117675
rect 12373 117663 12407 117675
rect 24624 115300 24696 119300
rect 24895 115333 25013 119267
rect 25284 115300 25344 119300
rect 25544 115300 25616 119300
rect 25815 115333 25933 119267
rect 26204 115300 26264 119300
rect 26464 115300 26536 119300
rect 26735 115333 26853 119267
rect 27124 115300 27184 119300
rect 27384 115300 27456 119300
rect 27655 115333 27773 119267
rect 28044 115300 28104 119300
rect 28304 115300 28376 119300
rect 28575 115333 28693 119267
rect 28964 115300 29024 119300
rect 29224 115300 29296 119300
rect 29495 115333 29613 119267
rect 29884 115300 29944 119300
rect 30144 115300 30216 119300
rect 30415 115333 30533 119267
rect 30804 115300 30864 119300
rect 31064 115300 31136 119300
rect 31335 115333 31453 119267
rect 31724 115300 31784 119300
rect 31984 115300 32056 119300
rect 32255 115333 32373 119267
rect 32644 115300 32704 119300
rect 59624 118764 59696 122764
rect 59895 118797 60013 122731
rect 60284 118764 60344 122764
rect 60544 118764 60616 122764
rect 60815 118797 60933 122731
rect 61204 118764 61264 122764
rect 61464 118764 61536 122764
rect 61735 118797 61853 122731
rect 62124 118764 62184 122764
rect 62384 118764 62456 122764
rect 62655 118797 62773 122731
rect 63044 118764 63104 122764
rect 63304 118764 63376 122764
rect 63575 118797 63693 122731
rect 63964 118764 64024 122764
rect 64224 118764 64296 122764
rect 64495 118797 64613 122731
rect 64884 118764 64944 122764
rect 65144 118764 65216 122764
rect 65415 118797 65533 122731
rect 65804 118764 65864 122764
rect 66064 118764 66136 122764
rect 66335 118797 66453 122731
rect 66724 118764 66784 122764
rect 66984 118764 67056 122764
rect 67255 118797 67373 122731
rect 67644 118764 67704 122764
rect 67904 118764 67976 122764
rect 68175 118797 68293 122731
rect 68564 118764 68624 122764
rect 68824 118764 68896 122764
rect 69095 118797 69213 122731
rect 69484 118764 69544 122764
rect 80176 119734 80248 123734
rect 80447 119767 80565 123701
rect 80836 119734 80896 123734
rect 81096 119734 81168 123734
rect 81367 119767 81485 123701
rect 81756 119734 81816 123734
rect 82016 119734 82088 123734
rect 82287 119767 82405 123701
rect 82676 119734 82736 123734
rect 82936 119734 83008 123734
rect 83207 119767 83325 123701
rect 83596 119734 83656 123734
rect 83856 119734 83928 123734
rect 84127 119767 84245 123701
rect 84516 119734 84576 123734
rect 84776 119734 84848 123734
rect 85047 119767 85165 123701
rect 85436 119734 85496 123734
rect 85696 119734 85768 123734
rect 85967 119767 86085 123701
rect 86356 119734 86416 123734
rect 86616 119734 86688 123734
rect 86887 119767 87005 123701
rect 87276 119734 87336 123734
rect 87536 119734 87608 123734
rect 87807 119767 87925 123701
rect 88196 119734 88256 123734
rect 88456 119734 88528 123734
rect 88727 119767 88845 123701
rect 89116 119734 89176 123734
rect 89376 119734 89448 123734
rect 89647 119767 89765 123701
rect 90036 119734 90096 123734
rect 100233 123696 100234 123720
rect 100314 123696 100315 123720
rect 101069 123696 101070 123720
rect 101150 123696 101151 123720
rect 101905 123696 101906 123720
rect 101986 123696 101987 123720
rect 102741 123696 102742 123720
rect 102822 123696 102823 123720
rect 103577 123696 103578 123720
rect 103658 123696 103659 123720
rect 104413 123696 104414 123720
rect 104494 123696 104495 123720
rect 105249 123696 105250 123720
rect 105330 123696 105331 123720
rect 106085 123696 106086 123720
rect 106166 123696 106167 123720
rect 106921 123696 106922 123720
rect 107002 123696 107003 123720
rect 107757 123696 107758 123720
rect 107838 123696 107839 123720
rect 108593 123696 108594 123720
rect 108674 123696 108675 123720
rect 109429 123696 109430 123720
rect 109510 123696 109511 123720
rect 110265 123696 110266 123720
rect 110346 123696 110347 123720
rect 100257 123672 100291 123684
rect 101093 123672 101127 123684
rect 101929 123672 101963 123684
rect 102765 123672 102799 123684
rect 103601 123672 103635 123684
rect 104437 123672 104471 123684
rect 105273 123672 105307 123684
rect 106109 123672 106143 123684
rect 106945 123672 106979 123684
rect 107781 123672 107815 123684
rect 108617 123672 108651 123684
rect 109453 123672 109487 123684
rect 110289 123672 110323 123684
rect 121219 123327 121429 123363
rect 133481 123327 133594 123363
rect 134043 123327 134325 123363
rect 120808 122327 120912 123327
rect 121008 122327 121080 123327
rect 121254 122327 121255 123327
rect 121296 122327 121352 123327
rect 121393 122327 121394 123327
rect 121654 122327 121714 123327
rect 121914 122327 121986 123327
rect 122216 122327 122272 123327
rect 122288 122327 122344 123327
rect 122646 122327 122706 123327
rect 122906 122327 122978 123327
rect 123208 122327 123264 123327
rect 123280 122327 123336 123327
rect 123638 122327 123698 123327
rect 123898 122327 123970 123327
rect 124200 122327 124256 123327
rect 124272 122327 124328 123327
rect 124630 122327 124690 123327
rect 124890 122327 124962 123327
rect 125192 122327 125248 123327
rect 125264 122327 125320 123327
rect 125622 122327 125682 123327
rect 125882 122327 125954 123327
rect 126184 122327 126240 123327
rect 126256 122327 126312 123327
rect 126614 122327 126674 123327
rect 126874 122327 126946 123327
rect 127176 122327 127232 123327
rect 127248 122327 127304 123327
rect 127606 122327 127666 123327
rect 127866 122327 127938 123327
rect 128168 122327 128224 123327
rect 128240 122327 128296 123327
rect 128598 122327 128658 123327
rect 128858 122327 128930 123327
rect 129160 122327 129216 123327
rect 129232 122327 129288 123327
rect 129590 122327 129650 123327
rect 129850 122327 129922 123327
rect 130152 122327 130208 123327
rect 130224 122327 130280 123327
rect 130582 122327 130642 123327
rect 130842 122327 130914 123327
rect 131144 122327 131200 123327
rect 131216 122327 131272 123327
rect 131574 122327 131634 123327
rect 131834 122327 131906 123327
rect 132136 122327 132192 123327
rect 132208 122327 132264 123327
rect 132566 122327 132626 123327
rect 132826 122327 132898 123327
rect 133128 122327 133184 123327
rect 133200 122327 133256 123327
rect 133481 122327 133517 123327
rect 133558 122327 133594 123327
rect 133818 122327 133890 123327
rect 134043 122327 134079 123327
rect 134120 122327 134176 123327
rect 134192 122327 134248 123327
rect 134289 122327 134325 123327
rect 134536 122327 134596 123327
rect 134632 122327 134736 123327
rect 140710 122462 140814 123462
rect 140910 122462 140982 123462
rect 121219 122291 121429 122327
rect 133481 122291 133594 122327
rect 134043 122291 134325 122327
rect 100233 121696 100234 121720
rect 100314 121696 100315 121720
rect 101069 121696 101070 121720
rect 101150 121696 101151 121720
rect 101905 121696 101906 121720
rect 101986 121696 101987 121720
rect 102741 121696 102742 121720
rect 102822 121696 102823 121720
rect 103577 121696 103578 121720
rect 103658 121696 103659 121720
rect 104413 121696 104414 121720
rect 104494 121696 104495 121720
rect 105249 121696 105250 121720
rect 105330 121696 105331 121720
rect 106085 121696 106086 121720
rect 106166 121696 106167 121720
rect 106921 121696 106922 121720
rect 107002 121696 107003 121720
rect 107757 121696 107758 121720
rect 107838 121696 107839 121720
rect 108593 121696 108594 121720
rect 108674 121696 108675 121720
rect 109429 121696 109430 121720
rect 109510 121696 109511 121720
rect 110265 121696 110266 121720
rect 110346 121696 110347 121720
rect 100257 121672 100291 121684
rect 101093 121672 101127 121684
rect 101929 121672 101963 121684
rect 102765 121672 102799 121684
rect 103601 121672 103635 121684
rect 104437 121672 104471 121684
rect 105273 121672 105307 121684
rect 106109 121672 106143 121684
rect 106945 121672 106979 121684
rect 107781 121672 107815 121684
rect 108617 121672 108651 121684
rect 109453 121672 109487 121684
rect 110289 121672 110323 121684
rect 140661 119964 140677 120030
rect 120631 119824 120647 119890
rect 122655 119824 122671 119890
rect 128822 119758 128838 119774
rect 101905 119696 101906 119720
rect 101986 119696 101987 119720
rect 102741 119696 102742 119720
rect 102822 119696 102823 119720
rect 103577 119696 103578 119720
rect 103658 119696 103659 119720
rect 104413 119696 104414 119720
rect 104494 119696 104495 119720
rect 105249 119696 105250 119720
rect 105330 119696 105331 119720
rect 106085 119696 106086 119720
rect 106166 119696 106167 119720
rect 106921 119696 106922 119720
rect 107002 119696 107003 119720
rect 107757 119696 107758 119720
rect 107838 119696 107839 119720
rect 108593 119696 108594 119720
rect 108674 119696 108675 119720
rect 109429 119696 109430 119720
rect 109510 119696 109511 119720
rect 110265 119696 110266 119720
rect 110346 119696 110347 119720
rect 101929 119672 101963 119684
rect 102765 119672 102799 119684
rect 103601 119672 103635 119684
rect 104437 119672 104471 119684
rect 105273 119672 105307 119684
rect 106109 119672 106143 119684
rect 106945 119672 106979 119684
rect 107781 119672 107815 119684
rect 108617 119672 108651 119684
rect 109453 119672 109487 119684
rect 110289 119672 110323 119684
rect 128720 119452 128838 119758
rect 128822 119436 128838 119452
rect 131010 119758 131026 119774
rect 131010 119452 131128 119758
rect 131010 119436 131026 119452
rect 42963 118532 42964 118556
rect 43044 118532 43045 118556
rect 43799 118532 43800 118556
rect 43880 118532 43881 118556
rect 44635 118532 44636 118556
rect 44716 118532 44717 118556
rect 45471 118532 45472 118556
rect 45552 118532 45553 118556
rect 46307 118532 46308 118556
rect 46388 118532 46389 118556
rect 47143 118532 47144 118556
rect 47224 118532 47225 118556
rect 47979 118532 47980 118556
rect 48060 118532 48061 118556
rect 48815 118532 48816 118556
rect 48896 118532 48897 118556
rect 49651 118532 49652 118556
rect 49732 118532 49733 118556
rect 50487 118532 50488 118556
rect 50568 118532 50569 118556
rect 51323 118532 51324 118556
rect 51404 118532 51405 118556
rect 42987 118508 43021 118520
rect 43823 118508 43857 118520
rect 44659 118508 44693 118520
rect 45495 118508 45529 118520
rect 46331 118508 46365 118520
rect 47167 118508 47201 118520
rect 48003 118508 48037 118520
rect 48839 118508 48873 118520
rect 49675 118508 49709 118520
rect 50511 118508 50545 118520
rect 51347 118508 51381 118520
rect 42963 116911 42964 116935
rect 43044 116911 43045 116935
rect 43799 116911 43800 116935
rect 43880 116911 43881 116935
rect 44635 116911 44636 116935
rect 44716 116911 44717 116935
rect 45471 116911 45472 116935
rect 45552 116911 45553 116935
rect 46307 116911 46308 116935
rect 46388 116911 46389 116935
rect 47143 116911 47144 116935
rect 47224 116911 47225 116935
rect 47979 116911 47980 116935
rect 48060 116911 48061 116935
rect 48815 116911 48816 116935
rect 48896 116911 48897 116935
rect 49651 116911 49652 116935
rect 49732 116911 49733 116935
rect 50487 116911 50488 116935
rect 50568 116911 50569 116935
rect 51323 116911 51324 116935
rect 51404 116911 51405 116935
rect 42987 116887 43021 116899
rect 43823 116887 43857 116899
rect 44659 116887 44693 116899
rect 45495 116887 45529 116899
rect 46331 116887 46365 116899
rect 47167 116887 47201 116899
rect 48003 116887 48037 116899
rect 48839 116887 48873 116899
rect 49675 116887 49709 116899
rect 50511 116887 50545 116899
rect 51347 116887 51381 116899
rect 24624 110700 24696 114700
rect 24895 110733 25013 114667
rect 25284 110700 25344 114700
rect 25544 110700 25616 114700
rect 25815 110733 25933 114667
rect 26204 110700 26264 114700
rect 26464 110700 26536 114700
rect 26735 110733 26853 114667
rect 27124 110700 27184 114700
rect 27384 110700 27456 114700
rect 27655 110733 27773 114667
rect 28044 110700 28104 114700
rect 28304 110700 28376 114700
rect 28575 110733 28693 114667
rect 28964 110700 29024 114700
rect 29224 110700 29296 114700
rect 29495 110733 29613 114667
rect 29884 110700 29944 114700
rect 30144 110700 30216 114700
rect 30415 110733 30533 114667
rect 30804 110700 30864 114700
rect 31064 110700 31136 114700
rect 31335 110733 31453 114667
rect 31724 110700 31784 114700
rect 31984 110700 32056 114700
rect 32255 110733 32373 114667
rect 32644 110700 32704 114700
rect 61464 114164 61536 118164
rect 61735 114197 61853 118131
rect 62124 114164 62184 118164
rect 62384 114164 62456 118164
rect 62655 114197 62773 118131
rect 63044 114164 63104 118164
rect 63304 114164 63376 118164
rect 63575 114197 63693 118131
rect 63964 114164 64024 118164
rect 64224 114164 64296 118164
rect 64495 114197 64613 118131
rect 64884 114164 64944 118164
rect 65144 114164 65216 118164
rect 65415 114197 65533 118131
rect 65804 114164 65864 118164
rect 66064 114164 66136 118164
rect 66335 114197 66453 118131
rect 66724 114164 66784 118164
rect 66984 114164 67056 118164
rect 67255 114197 67373 118131
rect 67644 114164 67704 118164
rect 67904 114164 67976 118164
rect 68175 114197 68293 118131
rect 68564 114164 68624 118164
rect 68824 114164 68896 118164
rect 69095 114197 69213 118131
rect 69484 114164 69544 118164
rect 82016 115134 82088 119134
rect 82287 115167 82405 119101
rect 82676 115134 82736 119134
rect 82936 115134 83008 119134
rect 83207 115167 83325 119101
rect 83596 115134 83656 119134
rect 83856 115134 83928 119134
rect 84127 115167 84245 119101
rect 84516 115134 84576 119134
rect 84776 115134 84848 119134
rect 85047 115167 85165 119101
rect 85436 115134 85496 119134
rect 85696 115134 85768 119134
rect 85967 115167 86085 119101
rect 86356 115134 86416 119134
rect 86616 115134 86688 119134
rect 86887 115167 87005 119101
rect 87276 115134 87336 119134
rect 87536 115134 87608 119134
rect 87807 115167 87925 119101
rect 88196 115134 88256 119134
rect 88456 115134 88528 119134
rect 88727 115167 88845 119101
rect 89116 115134 89176 119134
rect 89376 115134 89448 119134
rect 89647 115167 89765 119101
rect 90036 115134 90096 119134
rect 101905 118075 101906 118099
rect 101986 118075 101987 118099
rect 102741 118075 102742 118099
rect 102822 118075 102823 118099
rect 103577 118075 103578 118099
rect 103658 118075 103659 118099
rect 104413 118075 104414 118099
rect 104494 118075 104495 118099
rect 105249 118075 105250 118099
rect 105330 118075 105331 118099
rect 106085 118075 106086 118099
rect 106166 118075 106167 118099
rect 106921 118075 106922 118099
rect 107002 118075 107003 118099
rect 107757 118075 107758 118099
rect 107838 118075 107839 118099
rect 108593 118075 108594 118099
rect 108674 118075 108675 118099
rect 109429 118075 109430 118099
rect 109510 118075 109511 118099
rect 110265 118075 110266 118099
rect 110346 118075 110347 118099
rect 101929 118051 101963 118063
rect 102765 118051 102799 118063
rect 103601 118051 103635 118063
rect 104437 118051 104471 118063
rect 105273 118051 105307 118063
rect 106109 118051 106143 118063
rect 106945 118051 106979 118063
rect 107781 118051 107815 118063
rect 108617 118051 108651 118063
rect 109453 118051 109487 118063
rect 110289 118051 110323 118063
rect 120254 117573 120278 118362
rect 24624 106100 24696 110100
rect 24895 106133 25013 110067
rect 25284 106100 25344 110100
rect 25544 106100 25616 110100
rect 25815 106133 25933 110067
rect 26204 106100 26264 110100
rect 26464 106100 26536 110100
rect 26735 106133 26853 110067
rect 27124 106100 27184 110100
rect 27384 106100 27456 110100
rect 27655 106133 27773 110067
rect 28044 106100 28104 110100
rect 28304 106100 28376 110100
rect 28575 106133 28693 110067
rect 28964 106100 29024 110100
rect 29224 106100 29296 110100
rect 29495 106133 29613 110067
rect 29884 106100 29944 110100
rect 30144 106100 30216 110100
rect 30415 106133 30533 110067
rect 30804 106100 30864 110100
rect 31064 106100 31136 110100
rect 31335 106133 31453 110067
rect 31724 106100 31784 110100
rect 31984 106100 32056 110100
rect 32255 106133 32373 110067
rect 32644 106100 32704 110100
rect 61464 109564 61536 113564
rect 61735 109597 61853 113531
rect 62124 109564 62184 113564
rect 62384 109564 62456 113564
rect 62655 109597 62773 113531
rect 63044 109564 63104 113564
rect 63304 109564 63376 113564
rect 63575 109597 63693 113531
rect 63964 109564 64024 113564
rect 64224 109564 64296 113564
rect 64495 109597 64613 113531
rect 64884 109564 64944 113564
rect 65144 109564 65216 113564
rect 65415 109597 65533 113531
rect 65804 109564 65864 113564
rect 66064 109564 66136 113564
rect 66335 109597 66453 113531
rect 66724 109564 66784 113564
rect 66984 109564 67056 113564
rect 67255 109597 67373 113531
rect 67644 109564 67704 113564
rect 67904 109564 67976 113564
rect 68175 109597 68293 113531
rect 68564 109564 68624 113564
rect 68824 109564 68896 113564
rect 69095 109597 69213 113531
rect 69484 109564 69544 113564
rect 82016 110534 82088 114534
rect 82287 110567 82405 114501
rect 82676 110534 82736 114534
rect 82936 110534 83008 114534
rect 83207 110567 83325 114501
rect 83596 110534 83656 114534
rect 83856 110534 83928 114534
rect 84127 110567 84245 114501
rect 84516 110534 84576 114534
rect 84776 110534 84848 114534
rect 85047 110567 85165 114501
rect 85436 110534 85496 114534
rect 85696 110534 85768 114534
rect 85967 110567 86085 114501
rect 86356 110534 86416 114534
rect 86616 110534 86688 114534
rect 86887 110567 87005 114501
rect 87276 110534 87336 114534
rect 87536 110534 87608 114534
rect 87807 110567 87925 114501
rect 88196 110534 88256 114534
rect 88456 110534 88528 114534
rect 88727 110567 88845 114501
rect 89116 110534 89176 114534
rect 89376 110534 89448 114534
rect 89647 110567 89765 114501
rect 90036 110534 90096 114534
rect 120123 112827 120130 117570
rect 121583 116639 121695 116665
rect 121783 116639 121869 116665
rect 122575 116639 122687 116665
rect 122775 116639 122861 116665
rect 123567 116639 123679 116665
rect 123767 116639 123853 116665
rect 124559 116639 124671 116665
rect 124759 116639 124845 116665
rect 125551 116639 125663 116665
rect 125751 116639 125837 116665
rect 126543 116639 126655 116665
rect 126743 116639 126829 116665
rect 127535 116639 127647 116665
rect 127735 116639 127821 116665
rect 128527 116639 128639 116665
rect 128727 116639 128813 116665
rect 129519 116639 129631 116665
rect 129719 116639 129805 116665
rect 130511 116639 130623 116665
rect 130711 116639 130797 116665
rect 131503 116639 131615 116665
rect 131703 116639 131789 116665
rect 132495 116639 132607 116665
rect 132695 116639 132781 116665
rect 133487 116639 133599 116665
rect 133687 116639 133773 116665
rect 120918 115639 120968 116639
rect 121179 115639 121235 116639
rect 121251 115639 121307 116639
rect 121609 115675 121695 116639
rect 121809 115717 121810 116639
rect 121869 115717 122021 116639
rect 121809 115675 122021 115717
rect 121596 115651 121695 115675
rect 121800 115651 122021 115675
rect 121609 115639 121695 115651
rect 121809 115639 122021 115651
rect 122171 115639 122227 116639
rect 122243 115639 122299 116639
rect 122601 115675 122687 116639
rect 122801 115717 122802 116639
rect 122861 115717 123013 116639
rect 122801 115675 123013 115717
rect 122588 115651 122687 115675
rect 122792 115651 123013 115675
rect 122601 115639 122687 115651
rect 122801 115639 123013 115651
rect 123163 115639 123219 116639
rect 123235 115639 123291 116639
rect 123593 115675 123679 116639
rect 123793 115717 123794 116639
rect 123853 115717 124005 116639
rect 123793 115675 124005 115717
rect 123580 115651 123679 115675
rect 123784 115651 124005 115675
rect 123593 115639 123679 115651
rect 123793 115639 124005 115651
rect 124155 115639 124211 116639
rect 124227 115639 124283 116639
rect 124585 115675 124671 116639
rect 124785 115717 124786 116639
rect 124845 115717 124997 116639
rect 124785 115675 124997 115717
rect 124572 115651 124671 115675
rect 124776 115651 124997 115675
rect 124585 115639 124671 115651
rect 124785 115639 124997 115651
rect 125147 115639 125203 116639
rect 125219 115639 125275 116639
rect 125577 115675 125663 116639
rect 125777 115717 125778 116639
rect 125837 115717 125989 116639
rect 125777 115675 125989 115717
rect 125564 115651 125663 115675
rect 125768 115651 125989 115675
rect 125577 115639 125663 115651
rect 125777 115639 125989 115651
rect 126139 115639 126195 116639
rect 126211 115639 126267 116639
rect 126569 115675 126655 116639
rect 126769 115717 126770 116639
rect 126829 115717 126981 116639
rect 126769 115675 126981 115717
rect 126556 115651 126655 115675
rect 126760 115651 126981 115675
rect 126569 115639 126655 115651
rect 126769 115639 126981 115651
rect 127131 115639 127187 116639
rect 127203 115639 127259 116639
rect 127561 115675 127647 116639
rect 127761 115717 127762 116639
rect 127821 115717 127973 116639
rect 127761 115675 127973 115717
rect 127548 115651 127647 115675
rect 127752 115651 127973 115675
rect 127561 115639 127647 115651
rect 127761 115639 127973 115651
rect 128123 115639 128179 116639
rect 128195 115639 128251 116639
rect 128553 115675 128639 116639
rect 128753 115717 128754 116639
rect 128813 115717 128965 116639
rect 128753 115675 128965 115717
rect 128540 115651 128639 115675
rect 128744 115651 128965 115675
rect 128553 115639 128639 115651
rect 128753 115639 128965 115651
rect 129115 115639 129171 116639
rect 129187 115639 129243 116639
rect 129545 115675 129631 116639
rect 129745 115717 129746 116639
rect 129805 115717 129957 116639
rect 129745 115675 129957 115717
rect 129532 115651 129631 115675
rect 129736 115651 129957 115675
rect 129545 115639 129631 115651
rect 129745 115639 129957 115651
rect 130107 115639 130163 116639
rect 130179 115639 130235 116639
rect 130537 115675 130623 116639
rect 130737 115717 130738 116639
rect 130797 115717 130949 116639
rect 130737 115675 130949 115717
rect 130524 115651 130623 115675
rect 130728 115651 130949 115675
rect 130537 115639 130623 115651
rect 130737 115639 130949 115651
rect 131099 115639 131155 116639
rect 131171 115639 131227 116639
rect 131529 115675 131615 116639
rect 131729 115717 131730 116639
rect 131789 115717 131941 116639
rect 131729 115675 131941 115717
rect 131516 115651 131615 115675
rect 131720 115651 131941 115675
rect 131529 115639 131615 115651
rect 131729 115639 131941 115651
rect 132091 115639 132147 116639
rect 132163 115639 132219 116639
rect 132521 115675 132607 116639
rect 132721 115717 132722 116639
rect 132781 115717 132933 116639
rect 132721 115675 132933 115717
rect 132508 115651 132607 115675
rect 132712 115651 132933 115675
rect 132521 115639 132607 115651
rect 132721 115639 132933 115651
rect 133083 115639 133139 116639
rect 133155 115639 133211 116639
rect 133513 115675 133599 116639
rect 133713 115717 133714 116639
rect 133773 115717 133925 116639
rect 133713 115675 133925 115717
rect 133500 115651 133599 115675
rect 133704 115651 133925 115675
rect 133513 115639 133599 115651
rect 133713 115639 133925 115651
rect 134034 115639 134106 116639
rect 134172 115639 134189 116639
rect 134359 115639 134392 116639
rect 140248 116622 140282 116646
rect 134515 116447 134583 116473
rect 134515 116413 134549 116439
rect 121620 115627 121654 115639
rect 121824 115627 121858 115639
rect 122612 115627 122646 115639
rect 122816 115627 122850 115639
rect 123604 115627 123638 115639
rect 123808 115627 123842 115639
rect 124596 115627 124630 115639
rect 124800 115627 124834 115639
rect 125588 115627 125622 115639
rect 125792 115627 125826 115639
rect 126580 115627 126614 115639
rect 126784 115627 126818 115639
rect 127572 115627 127606 115639
rect 127776 115627 127810 115639
rect 128564 115627 128598 115639
rect 128768 115627 128802 115639
rect 129556 115627 129590 115639
rect 129760 115627 129794 115639
rect 130548 115627 130582 115639
rect 130752 115627 130786 115639
rect 131540 115627 131574 115639
rect 131744 115627 131778 115639
rect 132532 115627 132566 115639
rect 132736 115627 132770 115639
rect 133524 115627 133558 115639
rect 133728 115627 133762 115639
rect 121628 115113 121850 115191
rect 122620 115113 122842 115191
rect 123612 115113 123834 115191
rect 124604 115113 124826 115191
rect 125596 115113 125818 115191
rect 126588 115113 126810 115191
rect 127580 115113 127802 115191
rect 128572 115113 128794 115191
rect 129564 115113 129786 115191
rect 130556 115113 130778 115191
rect 131548 115113 131770 115191
rect 132540 115113 132762 115191
rect 133532 115113 133754 115191
rect 121583 115039 121695 115065
rect 121783 115039 121869 115065
rect 122575 115039 122687 115065
rect 122775 115039 122861 115065
rect 123567 115039 123679 115065
rect 123767 115039 123853 115065
rect 124559 115039 124671 115065
rect 124759 115039 124845 115065
rect 125551 115039 125663 115065
rect 125751 115039 125837 115065
rect 126543 115039 126655 115065
rect 126743 115039 126829 115065
rect 127535 115039 127647 115065
rect 127735 115039 127821 115065
rect 128527 115039 128639 115065
rect 128727 115039 128813 115065
rect 129519 115039 129631 115065
rect 129719 115039 129805 115065
rect 130511 115039 130623 115065
rect 130711 115039 130797 115065
rect 131503 115039 131615 115065
rect 131703 115039 131789 115065
rect 132495 115039 132607 115065
rect 132695 115039 132781 115065
rect 133487 115039 133599 115065
rect 133687 115039 133773 115065
rect 120918 114039 120968 115039
rect 121179 114039 121235 115039
rect 121251 114039 121307 115039
rect 121609 115027 121695 115039
rect 121809 115027 121810 115039
rect 121596 115003 121695 115027
rect 121800 115003 121810 115027
rect 121609 114039 121695 115003
rect 121809 114040 121810 115003
rect 121869 114040 122021 115039
rect 121809 114039 122021 114040
rect 122171 114039 122227 115039
rect 122243 114039 122299 115039
rect 122601 115027 122687 115039
rect 122801 115027 122802 115039
rect 122588 115003 122687 115027
rect 122792 115003 122802 115027
rect 122601 114039 122687 115003
rect 122801 114040 122802 115003
rect 122861 114040 123013 115039
rect 122801 114039 123013 114040
rect 123163 114039 123219 115039
rect 123235 114039 123291 115039
rect 123593 115027 123679 115039
rect 123793 115027 123794 115039
rect 123580 115003 123679 115027
rect 123784 115003 123794 115027
rect 123593 114039 123679 115003
rect 123793 114040 123794 115003
rect 123853 114040 124005 115039
rect 123793 114039 124005 114040
rect 124155 114039 124211 115039
rect 124227 114039 124283 115039
rect 124585 115027 124671 115039
rect 124785 115027 124786 115039
rect 124572 115003 124671 115027
rect 124776 115003 124786 115027
rect 124585 114039 124671 115003
rect 124785 114040 124786 115003
rect 124845 114040 124997 115039
rect 124785 114039 124997 114040
rect 125147 114039 125203 115039
rect 125219 114039 125275 115039
rect 125577 115027 125663 115039
rect 125777 115027 125778 115039
rect 125564 115003 125663 115027
rect 125768 115003 125778 115027
rect 125577 114039 125663 115003
rect 125777 114040 125778 115003
rect 125837 114040 125989 115039
rect 125777 114039 125989 114040
rect 126139 114039 126195 115039
rect 126211 114039 126267 115039
rect 126569 115027 126655 115039
rect 126769 115027 126770 115039
rect 126556 115003 126655 115027
rect 126760 115003 126770 115027
rect 126569 114039 126655 115003
rect 126769 114040 126770 115003
rect 126829 114040 126981 115039
rect 126769 114039 126981 114040
rect 127131 114039 127187 115039
rect 127203 114039 127259 115039
rect 127561 115027 127647 115039
rect 127761 115027 127762 115039
rect 127548 115003 127647 115027
rect 127752 115003 127762 115027
rect 127561 114039 127647 115003
rect 127761 114040 127762 115003
rect 127821 114040 127973 115039
rect 127761 114039 127973 114040
rect 128123 114039 128179 115039
rect 128195 114039 128251 115039
rect 128553 115027 128639 115039
rect 128753 115027 128754 115039
rect 128540 115003 128639 115027
rect 128744 115003 128754 115027
rect 128553 114039 128639 115003
rect 128753 114040 128754 115003
rect 128813 114040 128965 115039
rect 128753 114039 128965 114040
rect 129115 114039 129171 115039
rect 129187 114039 129243 115039
rect 129545 115027 129631 115039
rect 129745 115027 129746 115039
rect 129532 115003 129631 115027
rect 129736 115003 129746 115027
rect 129545 114039 129631 115003
rect 129745 114040 129746 115003
rect 129805 114040 129957 115039
rect 129745 114039 129957 114040
rect 130107 114039 130163 115039
rect 130179 114039 130235 115039
rect 130537 115027 130623 115039
rect 130737 115027 130738 115039
rect 130524 115003 130623 115027
rect 130728 115003 130738 115027
rect 130537 114039 130623 115003
rect 130737 114040 130738 115003
rect 130797 114040 130949 115039
rect 130737 114039 130949 114040
rect 131099 114039 131155 115039
rect 131171 114039 131227 115039
rect 131529 115027 131615 115039
rect 131729 115027 131730 115039
rect 131516 115003 131615 115027
rect 131720 115003 131730 115027
rect 131529 114039 131615 115003
rect 131729 114040 131730 115003
rect 131789 114040 131941 115039
rect 131729 114039 131941 114040
rect 132091 114039 132147 115039
rect 132163 114039 132219 115039
rect 132521 115027 132607 115039
rect 132721 115027 132722 115039
rect 132508 115003 132607 115027
rect 132712 115003 132722 115027
rect 132521 114039 132607 115003
rect 132721 114040 132722 115003
rect 132781 114040 132933 115039
rect 132721 114039 132933 114040
rect 133083 114039 133139 115039
rect 133155 114039 133211 115039
rect 133513 115027 133599 115039
rect 133713 115027 133714 115039
rect 133500 115003 133599 115027
rect 133704 115003 133714 115027
rect 133513 114039 133599 115003
rect 133713 114040 133714 115003
rect 133773 114040 133925 115039
rect 133713 114039 133925 114040
rect 134034 114039 134106 115039
rect 134172 114039 134189 115039
rect 134359 114039 134392 115039
rect 140288 112935 140316 116622
rect 140960 115574 141010 116574
rect 161216 116425 161255 124211
rect 161216 116369 161256 116425
rect 161270 116369 161280 124211
rect 161216 116333 161280 116369
rect 140960 113974 141010 114974
rect 140194 112931 140316 112935
rect 140194 112911 140288 112931
rect 140194 112905 140197 112911
rect 120123 112801 120278 112827
rect 120368 112801 127264 112837
rect 140224 112834 140227 112905
rect 120278 112770 120404 112801
rect 120425 112770 120459 112794
rect 120493 112770 120527 112794
rect 120561 112770 120595 112794
rect 120629 112770 120663 112794
rect 120697 112770 120731 112794
rect 120765 112770 120799 112794
rect 120833 112770 120867 112794
rect 120901 112770 120935 112794
rect 120969 112770 121003 112794
rect 121037 112770 121071 112794
rect 121105 112770 121139 112794
rect 121173 112770 121207 112794
rect 121241 112770 121275 112794
rect 121309 112770 121343 112794
rect 121377 112770 121411 112794
rect 121445 112770 121479 112794
rect 121513 112770 121547 112794
rect 121581 112770 121615 112794
rect 121649 112770 121683 112794
rect 121717 112770 121751 112794
rect 121785 112770 121819 112794
rect 121853 112770 121887 112794
rect 121921 112770 121955 112794
rect 121989 112770 122023 112794
rect 122057 112770 122091 112794
rect 122125 112770 122159 112794
rect 122193 112770 122227 112794
rect 122261 112770 122295 112794
rect 122329 112770 122363 112794
rect 122397 112770 122431 112794
rect 122465 112770 122499 112794
rect 122533 112770 122567 112794
rect 122601 112770 122635 112794
rect 122669 112770 122703 112794
rect 122737 112770 122771 112794
rect 122805 112770 122839 112794
rect 122873 112770 122907 112794
rect 122941 112770 122975 112794
rect 123009 112770 123043 112794
rect 123077 112770 123111 112794
rect 123145 112770 123179 112794
rect 123213 112770 123247 112794
rect 123281 112770 123315 112794
rect 123349 112770 123383 112794
rect 123417 112770 123451 112794
rect 123485 112770 123519 112794
rect 123553 112770 123587 112794
rect 123621 112770 123655 112794
rect 123689 112770 123723 112794
rect 123787 112770 123821 112794
rect 123855 112770 123889 112794
rect 123923 112770 123957 112794
rect 123991 112770 124025 112794
rect 124059 112770 124093 112794
rect 124127 112770 124161 112794
rect 124195 112770 124229 112794
rect 124263 112770 124297 112794
rect 124331 112770 124365 112794
rect 124399 112770 124433 112794
rect 124467 112770 124501 112794
rect 124535 112770 124569 112794
rect 124603 112770 124637 112794
rect 124671 112770 124705 112794
rect 124739 112770 124773 112794
rect 124807 112770 124841 112794
rect 124875 112770 124909 112794
rect 124943 112770 124977 112794
rect 125011 112770 125045 112794
rect 125079 112770 125113 112794
rect 125147 112770 125181 112794
rect 125215 112770 125249 112794
rect 125283 112770 125317 112794
rect 125351 112770 125385 112794
rect 125419 112770 125453 112794
rect 125487 112770 125521 112794
rect 125555 112770 125589 112794
rect 125623 112770 125657 112794
rect 125691 112770 125725 112794
rect 125759 112770 125793 112794
rect 125827 112770 125861 112794
rect 125895 112770 125929 112794
rect 125963 112770 125997 112794
rect 126031 112770 126065 112794
rect 126099 112770 126133 112794
rect 126167 112770 126201 112794
rect 126235 112770 126269 112794
rect 126303 112770 126337 112794
rect 126371 112770 126405 112794
rect 126439 112770 126473 112794
rect 126507 112770 126541 112794
rect 126575 112770 126609 112794
rect 126643 112770 126677 112794
rect 126711 112770 126745 112794
rect 126779 112770 126813 112794
rect 126847 112770 126881 112794
rect 126915 112770 126949 112794
rect 126983 112770 127017 112794
rect 127051 112770 127085 112794
rect 127119 112770 127153 112794
rect 127228 112770 127264 112801
rect 120368 112747 127264 112770
rect 120368 112734 120425 112747
rect 120459 112734 120493 112747
rect 120527 112734 120561 112747
rect 120595 112734 120629 112747
rect 120663 112734 120697 112747
rect 120731 112734 120765 112747
rect 120799 112734 120833 112747
rect 120867 112734 120901 112747
rect 120935 112734 120969 112747
rect 121003 112734 121037 112747
rect 121071 112734 121105 112747
rect 121139 112734 121173 112747
rect 121207 112734 121241 112747
rect 121275 112734 121309 112747
rect 121343 112734 121377 112747
rect 121411 112734 121445 112747
rect 121479 112734 121513 112747
rect 121547 112734 121581 112747
rect 121615 112734 121649 112747
rect 121683 112734 121717 112747
rect 121751 112734 121785 112747
rect 121819 112734 121853 112747
rect 121887 112734 121921 112747
rect 121955 112734 121989 112747
rect 122023 112734 122057 112747
rect 122091 112734 122125 112747
rect 122159 112734 122193 112747
rect 122227 112734 122261 112747
rect 122295 112734 122329 112747
rect 122363 112734 122397 112747
rect 122431 112734 122465 112747
rect 122499 112734 122533 112747
rect 122567 112734 122601 112747
rect 122635 112734 122669 112747
rect 122703 112734 122737 112747
rect 122771 112734 122805 112747
rect 122839 112734 122873 112747
rect 122907 112734 122941 112747
rect 122975 112734 123009 112747
rect 123043 112734 123077 112747
rect 123111 112734 123145 112747
rect 123179 112734 123213 112747
rect 123247 112734 123281 112747
rect 123315 112734 123349 112747
rect 123383 112734 123417 112747
rect 123451 112734 123485 112747
rect 123519 112734 123553 112747
rect 123587 112734 123621 112747
rect 123655 112734 123689 112747
rect 123723 112734 123787 112747
rect 123821 112734 123855 112747
rect 123889 112734 123923 112747
rect 123957 112734 123991 112747
rect 124025 112734 124059 112747
rect 124093 112734 124127 112747
rect 124161 112734 124195 112747
rect 124229 112734 124263 112747
rect 124297 112734 124331 112747
rect 124365 112734 124399 112747
rect 124433 112734 124467 112747
rect 124501 112734 124535 112747
rect 124569 112734 124603 112747
rect 124637 112734 124671 112747
rect 124705 112734 124739 112747
rect 124773 112734 124807 112747
rect 124841 112734 124875 112747
rect 124909 112734 124943 112747
rect 124977 112734 125011 112747
rect 125045 112734 125079 112747
rect 125113 112734 125147 112747
rect 125181 112734 125215 112747
rect 125249 112734 125283 112747
rect 125317 112734 125351 112747
rect 125385 112734 125419 112747
rect 125453 112734 125487 112747
rect 125521 112734 125555 112747
rect 125589 112734 125623 112747
rect 125657 112734 125691 112747
rect 125725 112734 125759 112747
rect 125793 112734 125827 112747
rect 125861 112734 125895 112747
rect 125929 112734 125963 112747
rect 125997 112734 126031 112747
rect 126065 112734 126099 112747
rect 126133 112734 126167 112747
rect 126201 112734 126235 112747
rect 126269 112734 126303 112747
rect 126337 112734 126371 112747
rect 126405 112734 126439 112747
rect 126473 112734 126507 112747
rect 126541 112734 126575 112747
rect 126609 112734 126643 112747
rect 126677 112734 126711 112747
rect 126745 112734 126779 112747
rect 126813 112734 126847 112747
rect 126881 112734 126915 112747
rect 126949 112734 126983 112747
rect 127017 112734 127051 112747
rect 127085 112734 127119 112747
rect 127153 112734 127264 112747
rect 121044 112423 122044 112473
rect 122174 112423 123574 112473
rect 123936 112423 125336 112473
rect 125466 112423 126866 112473
rect 121044 112267 122044 112395
rect 122174 112267 123574 112395
rect 123936 112267 125336 112395
rect 125466 112267 126866 112395
rect 121044 112111 122044 112239
rect 122174 112111 123574 112239
rect 123936 112111 125336 112239
rect 125466 112111 126866 112239
rect 121044 111955 122044 112083
rect 122174 111955 123574 112083
rect 123936 111955 125336 112083
rect 125466 111955 126866 112083
rect 128877 112031 129047 112337
rect 132165 112001 132181 112067
rect 134189 112001 134205 112067
rect 121044 111805 122044 111855
rect 122174 111805 123574 111855
rect 123936 111805 125336 111855
rect 125466 111805 126866 111855
rect 121202 111368 121236 111392
rect 121270 111368 121304 111392
rect 121338 111368 121372 111392
rect 121406 111368 121440 111392
rect 121474 111368 121508 111392
rect 121542 111368 121576 111392
rect 121610 111368 121644 111392
rect 121678 111368 121712 111392
rect 121746 111368 121780 111392
rect 121814 111368 121848 111392
rect 121882 111368 121916 111392
rect 121950 111368 121984 111392
rect 122018 111368 122052 111392
rect 122086 111368 122120 111392
rect 122154 111368 122188 111392
rect 122222 111368 122256 111392
rect 122290 111368 122324 111392
rect 122358 111368 122392 111392
rect 122426 111368 122460 111392
rect 122494 111368 122528 111392
rect 122562 111368 122596 111392
rect 122630 111368 122664 111392
rect 122698 111368 122732 111392
rect 122766 111368 122800 111392
rect 122834 111368 122868 111392
rect 122902 111368 122936 111392
rect 122970 111368 123004 111392
rect 123038 111368 123072 111392
rect 123106 111368 123140 111392
rect 123174 111368 123208 111392
rect 123242 111368 123276 111392
rect 123310 111368 123344 111392
rect 123378 111368 123412 111392
rect 123446 111368 123480 111392
rect 123514 111368 123548 111392
rect 123582 111368 123616 111392
rect 123650 111368 123684 111392
rect 123718 111368 123752 111392
rect 123786 111368 123820 111392
rect 123854 111368 123888 111392
rect 123922 111368 123956 111392
rect 123990 111368 124024 111392
rect 124058 111368 124092 111392
rect 124126 111368 124160 111392
rect 124194 111368 124228 111392
rect 124262 111368 124296 111392
rect 124330 111368 124364 111392
rect 124398 111368 124432 111392
rect 124466 111368 124500 111392
rect 124534 111368 124568 111392
rect 124602 111368 124636 111392
rect 124670 111368 124704 111392
rect 124738 111368 124772 111392
rect 124806 111368 124840 111392
rect 124874 111368 124908 111392
rect 124942 111368 124976 111392
rect 125010 111368 125044 111392
rect 125067 111343 125068 111368
rect 125026 111334 125068 111343
rect 121577 111004 124577 111054
rect 121577 110848 124577 110976
rect 125026 110932 125128 110956
rect 125026 110908 125050 110932
rect 125104 110908 125128 110932
rect 126509 110908 126543 110966
rect 126698 110932 126732 110966
rect 126770 110932 126804 110966
rect 126842 110932 126876 110966
rect 126914 110932 126948 110966
rect 126698 110908 126722 110932
rect 126924 110908 126948 110932
rect 127102 110932 127204 110956
rect 128332 110945 128356 110969
rect 128230 110932 128254 110935
rect 127102 110908 127126 110932
rect 127180 110908 127204 110932
rect 128308 110921 128332 110935
rect 128485 110932 128587 110956
rect 121577 110692 124577 110820
rect 121577 110536 124577 110664
rect 121577 110380 124577 110508
rect 121577 110224 124577 110352
rect 121577 110068 124577 110196
rect 1823 105308 1824 105332
rect 1904 105308 1905 105332
rect 2377 105308 2378 105332
rect 2458 105308 2459 105332
rect 2931 105308 2932 105332
rect 3012 105308 3013 105332
rect 3485 105308 3486 105332
rect 3566 105308 3567 105332
rect 4039 105308 4040 105332
rect 4120 105308 4121 105332
rect 4593 105308 4594 105332
rect 4674 105308 4675 105332
rect 5147 105308 5148 105332
rect 5228 105308 5229 105332
rect 5701 105308 5702 105332
rect 5782 105308 5783 105332
rect 6255 105308 6256 105332
rect 6336 105308 6337 105332
rect 6809 105308 6810 105332
rect 6890 105308 6891 105332
rect 7363 105308 7364 105332
rect 7444 105308 7445 105332
rect 7917 105308 7918 105332
rect 7998 105308 7999 105332
rect 8471 105308 8472 105332
rect 8552 105308 8553 105332
rect 9025 105308 9026 105332
rect 9106 105308 9107 105332
rect 9579 105308 9580 105332
rect 9660 105308 9661 105332
rect 10133 105308 10134 105332
rect 10214 105308 10215 105332
rect 10687 105308 10688 105332
rect 10768 105308 10769 105332
rect 11241 105308 11242 105332
rect 11322 105308 11323 105332
rect 11795 105308 11796 105332
rect 11876 105308 11877 105332
rect 12349 105308 12350 105332
rect 12430 105308 12431 105332
rect 1847 105284 1881 105296
rect 2401 105284 2435 105296
rect 2955 105284 2989 105296
rect 3509 105284 3543 105296
rect 4063 105284 4097 105296
rect 4617 105284 4651 105296
rect 5171 105284 5205 105296
rect 5725 105284 5759 105296
rect 6279 105284 6313 105296
rect 6833 105284 6867 105296
rect 7387 105284 7421 105296
rect 7941 105284 7975 105296
rect 8495 105284 8529 105296
rect 9049 105284 9083 105296
rect 9603 105284 9637 105296
rect 10157 105284 10191 105296
rect 10711 105284 10745 105296
rect 11265 105284 11299 105296
rect 11819 105284 11853 105296
rect 12373 105284 12407 105296
rect 1823 103308 1824 103332
rect 1904 103308 1905 103332
rect 2377 103308 2378 103332
rect 2458 103308 2459 103332
rect 2931 103308 2932 103332
rect 3012 103308 3013 103332
rect 3485 103308 3486 103332
rect 3566 103308 3567 103332
rect 4039 103308 4040 103332
rect 4120 103308 4121 103332
rect 4593 103308 4594 103332
rect 4674 103308 4675 103332
rect 5147 103308 5148 103332
rect 5228 103308 5229 103332
rect 5701 103308 5702 103332
rect 5782 103308 5783 103332
rect 6255 103308 6256 103332
rect 6336 103308 6337 103332
rect 6809 103308 6810 103332
rect 6890 103308 6891 103332
rect 7363 103308 7364 103332
rect 7444 103308 7445 103332
rect 7917 103308 7918 103332
rect 7998 103308 7999 103332
rect 8471 103308 8472 103332
rect 8552 103308 8553 103332
rect 9025 103308 9026 103332
rect 9106 103308 9107 103332
rect 9579 103308 9580 103332
rect 9660 103308 9661 103332
rect 10133 103308 10134 103332
rect 10214 103308 10215 103332
rect 10687 103308 10688 103332
rect 10768 103308 10769 103332
rect 11241 103308 11242 103332
rect 11322 103308 11323 103332
rect 11795 103308 11796 103332
rect 11876 103308 11877 103332
rect 12349 103308 12350 103332
rect 12430 103308 12431 103332
rect 1847 103284 1881 103296
rect 2401 103284 2435 103296
rect 2955 103284 2989 103296
rect 3509 103284 3543 103296
rect 4063 103284 4097 103296
rect 4617 103284 4651 103296
rect 5171 103284 5205 103296
rect 5725 103284 5759 103296
rect 6279 103284 6313 103296
rect 6833 103284 6867 103296
rect 7387 103284 7421 103296
rect 7941 103284 7975 103296
rect 8495 103284 8529 103296
rect 9049 103284 9083 103296
rect 9603 103284 9637 103296
rect 10157 103284 10191 103296
rect 10711 103284 10745 103296
rect 11265 103284 11299 103296
rect 11819 103284 11853 103296
rect 12373 103284 12407 103296
rect 22784 101500 22856 105500
rect 23055 101533 23173 105467
rect 23444 101500 23504 105500
rect 23704 101500 23776 105500
rect 23975 101533 24093 105467
rect 24364 101500 24424 105500
rect 24624 101500 24696 105500
rect 24895 101533 25013 105467
rect 25284 101500 25344 105500
rect 25544 101500 25616 105500
rect 25815 101533 25933 105467
rect 26204 101500 26264 105500
rect 26464 101500 26536 105500
rect 26735 101533 26853 105467
rect 27124 101500 27184 105500
rect 27384 101500 27456 105500
rect 27655 101533 27773 105467
rect 28044 101500 28104 105500
rect 28304 101500 28376 105500
rect 28575 101533 28693 105467
rect 28964 101500 29024 105500
rect 29224 101500 29296 105500
rect 29495 101533 29613 105467
rect 29884 101500 29944 105500
rect 30144 101500 30216 105500
rect 30415 101533 30533 105467
rect 30804 101500 30864 105500
rect 31064 101500 31136 105500
rect 31335 101533 31453 105467
rect 31724 101500 31784 105500
rect 31984 101500 32056 105500
rect 32255 101533 32373 105467
rect 32644 101500 32704 105500
rect 61464 104964 61536 108964
rect 61735 104997 61853 108931
rect 62124 104964 62184 108964
rect 62384 104964 62456 108964
rect 62655 104997 62773 108931
rect 63044 104964 63104 108964
rect 63304 104964 63376 108964
rect 63575 104997 63693 108931
rect 63964 104964 64024 108964
rect 64224 104964 64296 108964
rect 64495 104997 64613 108931
rect 64884 104964 64944 108964
rect 65144 104964 65216 108964
rect 65415 104997 65533 108931
rect 65804 104964 65864 108964
rect 66064 104964 66136 108964
rect 66335 104997 66453 108931
rect 66724 104964 66784 108964
rect 66984 104964 67056 108964
rect 67255 104997 67373 108931
rect 67644 104964 67704 108964
rect 67904 104964 67976 108964
rect 68175 104997 68293 108931
rect 68564 104964 68624 108964
rect 68824 104964 68896 108964
rect 69095 104997 69213 108931
rect 69484 104964 69544 108964
rect 82016 105934 82088 109934
rect 82287 105967 82405 109901
rect 82676 105934 82736 109934
rect 82936 105934 83008 109934
rect 83207 105967 83325 109901
rect 83596 105934 83656 109934
rect 83856 105934 83928 109934
rect 84127 105967 84245 109901
rect 84516 105934 84576 109934
rect 84776 105934 84848 109934
rect 85047 105967 85165 109901
rect 85436 105934 85496 109934
rect 85696 105934 85768 109934
rect 85967 105967 86085 109901
rect 86356 105934 86416 109934
rect 86616 105934 86688 109934
rect 86887 105967 87005 109901
rect 87276 105934 87336 109934
rect 87536 105934 87608 109934
rect 87807 105967 87925 109901
rect 88196 105934 88256 109934
rect 88456 105934 88528 109934
rect 88727 105967 88845 109901
rect 89116 105934 89176 109934
rect 89376 105934 89448 109934
rect 89647 105967 89765 109901
rect 90036 105934 90096 109934
rect 121577 109918 124577 109968
rect 125414 109504 125457 110904
rect 125564 109504 125692 110904
rect 125727 109504 125855 110904
rect 125890 109504 126018 110904
rect 126053 109504 126181 110904
rect 126216 109504 126344 110904
rect 126379 109504 126422 110904
rect 127291 109504 127341 110904
rect 127448 109504 127576 110904
rect 127611 109504 127739 110904
rect 127774 109504 127902 110904
rect 127937 109504 128065 110904
rect 128100 109504 128143 110904
rect 128206 110887 128230 110911
rect 128332 110887 128356 110911
rect 128485 110908 128509 110932
rect 128563 110908 128587 110932
rect 122070 109105 122240 109411
rect 122870 109105 123040 109411
rect 123670 109105 123840 109411
rect 122070 108605 122240 108911
rect 122870 108605 123040 108911
rect 123670 108605 123840 108911
rect 119527 107145 119577 107745
rect 119677 107145 119805 107745
rect 119833 107145 119961 107745
rect 119989 107145 120045 107745
rect 120145 107145 120273 107745
rect 120301 107145 120429 107745
rect 120457 107145 120507 107745
rect 120587 107145 120637 107745
rect 120737 107145 120787 107745
rect 121225 107144 121275 107744
rect 121375 107144 121503 107744
rect 121531 107144 121659 107744
rect 121687 107144 121743 107744
rect 121843 107144 121971 107744
rect 121999 107144 122127 107744
rect 122155 107144 122205 107744
rect 122285 107144 122335 107744
rect 122435 107144 122485 107744
rect 122607 107144 122657 107744
rect 122757 107144 122807 107744
rect 122887 107144 122937 107744
rect 123037 107144 123165 107744
rect 123193 107144 123321 107744
rect 123349 107144 123405 107744
rect 123505 107144 123633 107744
rect 123661 107144 123789 107744
rect 123817 107144 123867 107744
rect 125414 107232 125457 108632
rect 125564 107232 125692 108632
rect 125727 107232 125855 108632
rect 125890 107232 126018 108632
rect 126053 107232 126181 108632
rect 126216 107232 126344 108632
rect 126379 107232 126422 108632
rect 125026 107204 125128 107228
rect 125104 107180 125128 107204
rect 126509 107180 126543 107238
rect 126698 107204 126732 107238
rect 126770 107204 126804 107238
rect 126842 107204 126876 107238
rect 126914 107204 126948 107238
rect 127291 107232 127341 108632
rect 127448 107232 127576 108632
rect 127611 107232 127739 108632
rect 127774 107232 127902 108632
rect 127937 107232 128065 108632
rect 128100 107232 128143 108632
rect 126698 107180 126722 107204
rect 126924 107180 126948 107204
rect 127102 107204 127204 107228
rect 128206 107225 128230 107249
rect 128332 107225 128356 107249
rect 127102 107180 127126 107204
rect 127180 107180 127204 107204
rect 128230 107201 128254 107204
rect 128308 107201 128332 107215
rect 128485 107204 128587 107228
rect 128332 107167 128356 107191
rect 128485 107180 128509 107204
rect 128563 107180 128587 107204
rect 128763 106764 129299 111372
rect 131734 111064 131825 111166
rect 132058 111131 132072 111155
rect 132024 111107 132048 111131
rect 132082 111107 132106 111131
rect 135278 111057 135312 111077
rect 131681 110944 131705 110968
rect 131739 110944 131763 110968
rect 132215 110962 132249 110966
rect 132283 110962 132317 110966
rect 132351 110962 132385 110966
rect 132419 110962 132453 110966
rect 132487 110962 132521 110966
rect 132555 110962 132589 110966
rect 132623 110962 132657 110966
rect 132691 110962 132725 110966
rect 132759 110962 132793 110966
rect 132827 110962 132861 110966
rect 132895 110962 132929 110966
rect 132963 110962 132997 110966
rect 133031 110962 133065 110966
rect 133099 110962 133133 110966
rect 133167 110962 133201 110966
rect 133235 110962 133269 110966
rect 133303 110962 133337 110966
rect 133371 110962 133405 110966
rect 133439 110962 133473 110966
rect 133507 110962 133541 110966
rect 133575 110962 133609 110966
rect 133643 110962 133677 110966
rect 133711 110962 133745 110966
rect 133779 110962 133813 110966
rect 133847 110962 133881 110966
rect 133915 110962 133949 110966
rect 133983 110962 134017 110966
rect 134051 110962 134085 110966
rect 134119 110962 134153 110966
rect 134187 110962 134221 110966
rect 134255 110962 134289 110966
rect 134323 110962 134357 110966
rect 134391 110962 134425 110966
rect 134459 110962 134493 110966
rect 134527 110962 134561 110966
rect 134595 110962 134629 110966
rect 134663 110962 134697 110966
rect 134731 110962 134765 110966
rect 134799 110962 134833 110966
rect 134867 110962 134901 110966
rect 134935 110962 134969 110966
rect 132147 110944 135047 110962
rect 132215 110940 132249 110944
rect 132283 110940 132317 110944
rect 132351 110940 132385 110944
rect 132419 110940 132453 110944
rect 132487 110940 132521 110944
rect 132555 110940 132589 110944
rect 132623 110940 132657 110944
rect 132691 110940 132725 110944
rect 132759 110940 132793 110944
rect 132827 110940 132861 110944
rect 132895 110940 132929 110944
rect 132963 110940 132997 110944
rect 133031 110940 133065 110944
rect 133099 110940 133133 110944
rect 133167 110940 133201 110944
rect 133235 110940 133269 110944
rect 133303 110940 133337 110944
rect 133371 110940 133405 110944
rect 133439 110940 133473 110944
rect 133507 110940 133541 110944
rect 133575 110940 133609 110944
rect 133643 110940 133677 110944
rect 133711 110940 133745 110944
rect 133779 110940 133813 110944
rect 133847 110940 133881 110944
rect 133915 110940 133949 110944
rect 133983 110940 134017 110944
rect 134051 110940 134085 110944
rect 134119 110940 134153 110944
rect 134187 110940 134221 110944
rect 134255 110940 134289 110944
rect 134323 110940 134357 110944
rect 134391 110940 134425 110944
rect 134459 110940 134493 110944
rect 134527 110940 134561 110944
rect 134595 110940 134629 110944
rect 134663 110940 134697 110944
rect 134731 110940 134765 110944
rect 134799 110940 134833 110944
rect 134867 110940 134901 110944
rect 134935 110940 134969 110944
rect 135186 110941 135210 110965
rect 131705 110920 131739 110934
rect 132151 110932 135043 110940
rect 132191 110920 134993 110932
rect 135210 110917 135234 110932
rect 135278 110921 135312 110956
rect 129333 109504 129461 110904
rect 129496 109504 129624 110904
rect 129659 109504 129787 110904
rect 129822 109504 129950 110904
rect 129985 109504 130113 110904
rect 130148 109504 130276 110904
rect 130311 109504 130354 110904
rect 130447 109504 130490 110904
rect 130597 109504 130725 110904
rect 130760 109504 130888 110904
rect 130923 109504 131051 110904
rect 131086 109504 131214 110904
rect 131249 109504 131377 110904
rect 131412 109504 131540 110904
rect 131575 109504 131625 110904
rect 131681 110886 131705 110910
rect 131739 110886 131763 110910
rect 135288 110908 135312 110921
rect 131892 109119 131994 110683
rect 132261 109436 132311 110836
rect 132418 109436 132546 110836
rect 132581 109436 132709 110836
rect 132744 109436 132872 110836
rect 132907 109436 133035 110836
rect 133070 109436 133198 110836
rect 133233 109436 133361 110836
rect 133396 109436 133439 110836
rect 133532 109436 133575 110836
rect 133682 109436 133810 110836
rect 133845 109436 133973 110836
rect 134008 109436 134136 110836
rect 134171 109436 134299 110836
rect 134334 109436 134462 110836
rect 134497 109436 134625 110836
rect 134660 109436 134788 110836
rect 134823 109436 134866 110836
rect 140951 109684 140967 109750
rect 131926 109095 131960 109119
rect 131926 109017 131960 109041
rect 129333 107232 129461 108632
rect 129496 107232 129624 108632
rect 129659 107232 129787 108632
rect 129822 107232 129950 108632
rect 129985 107232 130113 108632
rect 130148 107232 130276 108632
rect 130311 107232 130354 108632
rect 130447 107232 130490 108632
rect 130597 107232 130725 108632
rect 130760 107232 130888 108632
rect 130923 107232 131051 108632
rect 131086 107232 131214 108632
rect 131249 107232 131377 108632
rect 131412 107232 131540 108632
rect 131575 107232 131625 108632
rect 131892 107453 131994 109017
rect 132261 107300 132311 108700
rect 132418 107300 132546 108700
rect 132581 107300 132709 108700
rect 132744 107300 132872 108700
rect 132907 107300 133035 108700
rect 133070 107300 133198 108700
rect 133233 107300 133361 108700
rect 133396 107300 133439 108700
rect 133532 107300 133575 108700
rect 133682 107300 133810 108700
rect 133845 107300 133973 108700
rect 134008 107300 134136 108700
rect 134171 107300 134299 108700
rect 134334 107300 134462 108700
rect 134497 107300 134625 108700
rect 134660 107300 134788 108700
rect 134823 107300 134866 108700
rect 131681 107226 131705 107250
rect 131739 107226 131763 107250
rect 132215 107234 132249 107238
rect 132283 107234 132317 107238
rect 132351 107234 132385 107238
rect 132419 107234 132453 107238
rect 132487 107234 132521 107238
rect 132555 107234 132589 107238
rect 132623 107234 132657 107238
rect 132691 107234 132725 107238
rect 132759 107234 132793 107238
rect 132827 107234 132861 107238
rect 132895 107234 132929 107238
rect 132963 107234 132997 107238
rect 133031 107234 133065 107238
rect 133099 107234 133133 107238
rect 133167 107234 133201 107238
rect 133235 107234 133269 107238
rect 133303 107234 133337 107238
rect 133371 107234 133405 107238
rect 133439 107234 133473 107238
rect 133507 107234 133541 107238
rect 133575 107234 133609 107238
rect 133643 107234 133677 107238
rect 133711 107234 133745 107238
rect 133779 107234 133813 107238
rect 133847 107234 133881 107238
rect 133915 107234 133949 107238
rect 133983 107234 134017 107238
rect 134051 107234 134085 107238
rect 134119 107234 134153 107238
rect 134187 107234 134221 107238
rect 134255 107234 134289 107238
rect 134323 107234 134357 107238
rect 134391 107234 134425 107238
rect 134459 107234 134493 107238
rect 134527 107234 134561 107238
rect 134595 107234 134629 107238
rect 134663 107234 134697 107238
rect 134731 107234 134765 107238
rect 134799 107234 134833 107238
rect 134867 107234 134901 107238
rect 134935 107234 134969 107238
rect 132181 107226 135013 107234
rect 135244 107229 135312 107249
rect 132215 107222 132249 107226
rect 132283 107222 132317 107226
rect 132351 107222 132385 107226
rect 132419 107222 132453 107226
rect 132487 107222 132521 107226
rect 132555 107222 132589 107226
rect 132623 107222 132657 107226
rect 132691 107222 132725 107226
rect 132759 107222 132793 107226
rect 132827 107222 132861 107226
rect 132895 107222 132929 107226
rect 132963 107222 132997 107226
rect 133031 107222 133065 107226
rect 133099 107222 133133 107226
rect 133167 107222 133201 107226
rect 133235 107222 133269 107226
rect 133303 107222 133337 107226
rect 133371 107222 133405 107226
rect 133439 107222 133473 107226
rect 133507 107222 133541 107226
rect 133575 107222 133609 107226
rect 133643 107222 133677 107226
rect 133711 107222 133745 107226
rect 133779 107222 133813 107226
rect 133847 107222 133881 107226
rect 133915 107222 133949 107226
rect 133983 107222 134017 107226
rect 134051 107222 134085 107226
rect 134119 107222 134153 107226
rect 134187 107222 134221 107226
rect 134255 107222 134289 107226
rect 134323 107222 134357 107226
rect 134391 107222 134425 107226
rect 134459 107222 134493 107226
rect 134527 107222 134561 107226
rect 134595 107222 134629 107226
rect 134663 107222 134697 107226
rect 134731 107222 134765 107226
rect 134799 107222 134833 107226
rect 134867 107222 134901 107226
rect 134935 107222 134969 107226
rect 131705 107202 131739 107216
rect 132147 107204 135047 107222
rect 135210 107204 135234 107219
rect 135278 107204 135312 107229
rect 132191 107202 134993 107204
rect 131681 107168 131705 107192
rect 131739 107168 131763 107192
rect 135186 107171 135210 107195
rect 135288 107180 135312 107204
rect 135244 107093 135312 107113
rect 131734 106970 131825 107072
rect 132024 107005 132048 107029
rect 132082 107005 132106 107029
rect 132058 106981 132072 107005
rect 99739 105696 99740 105720
rect 99820 105696 99821 105720
rect 100293 105696 100294 105720
rect 100374 105696 100375 105720
rect 100847 105696 100848 105720
rect 100928 105696 100929 105720
rect 101401 105696 101402 105720
rect 101482 105696 101483 105720
rect 101955 105696 101956 105720
rect 102036 105696 102037 105720
rect 102509 105696 102510 105720
rect 102590 105696 102591 105720
rect 103063 105696 103064 105720
rect 103144 105696 103145 105720
rect 103617 105696 103618 105720
rect 103698 105696 103699 105720
rect 104171 105696 104172 105720
rect 104252 105696 104253 105720
rect 104725 105696 104726 105720
rect 104806 105696 104807 105720
rect 105279 105696 105280 105720
rect 105360 105696 105361 105720
rect 105833 105696 105834 105720
rect 105914 105696 105915 105720
rect 106387 105696 106388 105720
rect 106468 105696 106469 105720
rect 106941 105696 106942 105720
rect 107022 105696 107023 105720
rect 107495 105696 107496 105720
rect 107576 105696 107577 105720
rect 108049 105696 108050 105720
rect 108130 105696 108131 105720
rect 108603 105696 108604 105720
rect 108684 105696 108685 105720
rect 109157 105696 109158 105720
rect 109238 105696 109239 105720
rect 109711 105696 109712 105720
rect 109792 105696 109793 105720
rect 110265 105696 110266 105720
rect 110346 105696 110347 105720
rect 99763 105672 99797 105684
rect 100317 105672 100351 105684
rect 100871 105672 100905 105684
rect 101425 105672 101459 105684
rect 101979 105672 102013 105684
rect 102533 105672 102567 105684
rect 103087 105672 103121 105684
rect 103641 105672 103675 105684
rect 104195 105672 104229 105684
rect 104749 105672 104783 105684
rect 105303 105672 105337 105684
rect 105857 105672 105891 105684
rect 106411 105672 106445 105684
rect 106965 105672 106999 105684
rect 107519 105672 107553 105684
rect 108073 105672 108107 105684
rect 108627 105672 108661 105684
rect 109181 105672 109215 105684
rect 109735 105672 109769 105684
rect 110289 105672 110323 105684
rect 121923 105627 121973 105827
rect 122073 105627 122129 105827
rect 122229 105627 122279 105827
rect 122629 105627 122679 105827
rect 122779 105627 122835 105827
rect 122935 105627 122985 105827
rect 123049 105627 123060 105827
rect 129913 105381 129963 106381
rect 130063 105381 130119 106381
rect 130219 105381 130275 106381
rect 130375 105381 130431 106381
rect 130531 105924 130581 106381
rect 130995 105924 131045 106381
rect 130531 105840 130584 105924
rect 130992 105840 131045 105924
rect 130531 105591 130581 105840
rect 130995 105591 131045 105840
rect 130531 105507 130584 105591
rect 130992 105507 131045 105591
rect 130531 105381 130581 105507
rect 130995 105381 131045 105507
rect 131145 105381 131201 106381
rect 131301 105381 131357 106381
rect 131457 105381 131513 106381
rect 131613 105381 131663 106381
rect 133848 105992 133898 106592
rect 133998 105992 134048 106592
rect 134120 105992 134170 106592
rect 134270 105992 134320 106592
rect 134396 105992 134446 106592
rect 134546 105992 134596 106592
rect 134668 105992 134718 106592
rect 134818 105992 134868 106592
rect 132804 105669 133110 105839
rect 40797 104532 40798 104556
rect 40878 104532 40879 104556
rect 41351 104532 41352 104556
rect 41432 104532 41433 104556
rect 41905 104532 41906 104556
rect 41986 104532 41987 104556
rect 42459 104532 42460 104556
rect 42540 104532 42541 104556
rect 43013 104532 43014 104556
rect 43094 104532 43095 104556
rect 43567 104532 43568 104556
rect 43648 104532 43649 104556
rect 44121 104532 44122 104556
rect 44202 104532 44203 104556
rect 44675 104532 44676 104556
rect 44756 104532 44757 104556
rect 45229 104532 45230 104556
rect 45310 104532 45311 104556
rect 45783 104532 45784 104556
rect 45864 104532 45865 104556
rect 46337 104532 46338 104556
rect 46418 104532 46419 104556
rect 46891 104532 46892 104556
rect 46972 104532 46973 104556
rect 47445 104532 47446 104556
rect 47526 104532 47527 104556
rect 47999 104532 48000 104556
rect 48080 104532 48081 104556
rect 48553 104532 48554 104556
rect 48634 104532 48635 104556
rect 49107 104532 49108 104556
rect 49188 104532 49189 104556
rect 49661 104532 49662 104556
rect 49742 104532 49743 104556
rect 50215 104532 50216 104556
rect 50296 104532 50297 104556
rect 50769 104532 50770 104556
rect 50850 104532 50851 104556
rect 51323 104532 51324 104556
rect 51404 104532 51405 104556
rect 40821 104508 40855 104520
rect 41375 104508 41409 104520
rect 41929 104508 41963 104520
rect 42483 104508 42517 104520
rect 43037 104508 43071 104520
rect 43591 104508 43625 104520
rect 44145 104508 44179 104520
rect 44699 104508 44733 104520
rect 45253 104508 45287 104520
rect 45807 104508 45841 104520
rect 46361 104508 46395 104520
rect 46915 104508 46949 104520
rect 47469 104508 47503 104520
rect 48023 104508 48057 104520
rect 48577 104508 48611 104520
rect 49131 104508 49165 104520
rect 49685 104508 49719 104520
rect 50239 104508 50273 104520
rect 50793 104508 50827 104520
rect 51347 104508 51381 104520
rect 40797 102532 40798 102556
rect 40878 102532 40879 102556
rect 41351 102532 41352 102556
rect 41432 102532 41433 102556
rect 41905 102532 41906 102556
rect 41986 102532 41987 102556
rect 42459 102532 42460 102556
rect 42540 102532 42541 102556
rect 43013 102532 43014 102556
rect 43094 102532 43095 102556
rect 43567 102532 43568 102556
rect 43648 102532 43649 102556
rect 44121 102532 44122 102556
rect 44202 102532 44203 102556
rect 44675 102532 44676 102556
rect 44756 102532 44757 102556
rect 45229 102532 45230 102556
rect 45310 102532 45311 102556
rect 45783 102532 45784 102556
rect 45864 102532 45865 102556
rect 46337 102532 46338 102556
rect 46418 102532 46419 102556
rect 46891 102532 46892 102556
rect 46972 102532 46973 102556
rect 47445 102532 47446 102556
rect 47526 102532 47527 102556
rect 47999 102532 48000 102556
rect 48080 102532 48081 102556
rect 48553 102532 48554 102556
rect 48634 102532 48635 102556
rect 49107 102532 49108 102556
rect 49188 102532 49189 102556
rect 49661 102532 49662 102556
rect 49742 102532 49743 102556
rect 50215 102532 50216 102556
rect 50296 102532 50297 102556
rect 50769 102532 50770 102556
rect 50850 102532 50851 102556
rect 51323 102532 51324 102556
rect 51404 102532 51405 102556
rect 40821 102508 40855 102520
rect 41375 102508 41409 102520
rect 41929 102508 41963 102520
rect 42483 102508 42517 102520
rect 43037 102508 43071 102520
rect 43591 102508 43625 102520
rect 44145 102508 44179 102520
rect 44699 102508 44733 102520
rect 45253 102508 45287 102520
rect 45807 102508 45841 102520
rect 46361 102508 46395 102520
rect 46915 102508 46949 102520
rect 47469 102508 47503 102520
rect 48023 102508 48057 102520
rect 48577 102508 48611 102520
rect 49131 102508 49165 102520
rect 49685 102508 49719 102520
rect 50239 102508 50273 102520
rect 50793 102508 50827 102520
rect 51347 102508 51381 102520
rect 1823 101308 1824 101332
rect 1904 101308 1905 101332
rect 2377 101308 2378 101332
rect 2458 101308 2459 101332
rect 2931 101308 2932 101332
rect 3012 101308 3013 101332
rect 3485 101308 3486 101332
rect 3566 101308 3567 101332
rect 4039 101308 4040 101332
rect 4120 101308 4121 101332
rect 4593 101308 4594 101332
rect 4674 101308 4675 101332
rect 5147 101308 5148 101332
rect 5228 101308 5229 101332
rect 5701 101308 5702 101332
rect 5782 101308 5783 101332
rect 6255 101308 6256 101332
rect 6336 101308 6337 101332
rect 6809 101308 6810 101332
rect 6890 101308 6891 101332
rect 7363 101308 7364 101332
rect 7444 101308 7445 101332
rect 7917 101308 7918 101332
rect 7998 101308 7999 101332
rect 8471 101308 8472 101332
rect 8552 101308 8553 101332
rect 9025 101308 9026 101332
rect 9106 101308 9107 101332
rect 9579 101308 9580 101332
rect 9660 101308 9661 101332
rect 10133 101308 10134 101332
rect 10214 101308 10215 101332
rect 10687 101308 10688 101332
rect 10768 101308 10769 101332
rect 11241 101308 11242 101332
rect 11322 101308 11323 101332
rect 11795 101308 11796 101332
rect 11876 101308 11877 101332
rect 12349 101308 12350 101332
rect 12430 101308 12431 101332
rect 1847 101284 1881 101296
rect 2401 101284 2435 101296
rect 2955 101284 2989 101296
rect 3509 101284 3543 101296
rect 4063 101284 4097 101296
rect 4617 101284 4651 101296
rect 5171 101284 5205 101296
rect 5725 101284 5759 101296
rect 6279 101284 6313 101296
rect 6833 101284 6867 101296
rect 7387 101284 7421 101296
rect 7941 101284 7975 101296
rect 8495 101284 8529 101296
rect 9049 101284 9083 101296
rect 9603 101284 9637 101296
rect 10157 101284 10191 101296
rect 10711 101284 10745 101296
rect 11265 101284 11299 101296
rect 11819 101284 11853 101296
rect 12373 101284 12407 101296
rect 40797 100532 40798 100556
rect 40878 100532 40879 100556
rect 41351 100532 41352 100556
rect 41432 100532 41433 100556
rect 41905 100532 41906 100556
rect 41986 100532 41987 100556
rect 42459 100532 42460 100556
rect 42540 100532 42541 100556
rect 43013 100532 43014 100556
rect 43094 100532 43095 100556
rect 43567 100532 43568 100556
rect 43648 100532 43649 100556
rect 44121 100532 44122 100556
rect 44202 100532 44203 100556
rect 44675 100532 44676 100556
rect 44756 100532 44757 100556
rect 45229 100532 45230 100556
rect 45310 100532 45311 100556
rect 45783 100532 45784 100556
rect 45864 100532 45865 100556
rect 46337 100532 46338 100556
rect 46418 100532 46419 100556
rect 46891 100532 46892 100556
rect 46972 100532 46973 100556
rect 47445 100532 47446 100556
rect 47526 100532 47527 100556
rect 47999 100532 48000 100556
rect 48080 100532 48081 100556
rect 48553 100532 48554 100556
rect 48634 100532 48635 100556
rect 49107 100532 49108 100556
rect 49188 100532 49189 100556
rect 49661 100532 49662 100556
rect 49742 100532 49743 100556
rect 50215 100532 50216 100556
rect 50296 100532 50297 100556
rect 50769 100532 50770 100556
rect 50850 100532 50851 100556
rect 51323 100532 51324 100556
rect 51404 100532 51405 100556
rect 40821 100508 40855 100520
rect 41375 100508 41409 100520
rect 41929 100508 41963 100520
rect 42483 100508 42517 100520
rect 43037 100508 43071 100520
rect 43591 100508 43625 100520
rect 44145 100508 44179 100520
rect 44699 100508 44733 100520
rect 45253 100508 45287 100520
rect 45807 100508 45841 100520
rect 46361 100508 46395 100520
rect 46915 100508 46949 100520
rect 47469 100508 47503 100520
rect 48023 100508 48057 100520
rect 48577 100508 48611 100520
rect 49131 100508 49165 100520
rect 49685 100508 49719 100520
rect 50239 100508 50273 100520
rect 50793 100508 50827 100520
rect 51347 100508 51381 100520
rect 59624 100364 59696 104364
rect 59895 100397 60013 104331
rect 60284 100364 60344 104364
rect 60544 100364 60616 104364
rect 60815 100397 60933 104331
rect 61204 100364 61264 104364
rect 61464 100364 61536 104364
rect 61735 100397 61853 104331
rect 62124 100364 62184 104364
rect 62384 100364 62456 104364
rect 62655 100397 62773 104331
rect 63044 100364 63104 104364
rect 63304 100364 63376 104364
rect 63575 100397 63693 104331
rect 63964 100364 64024 104364
rect 64224 100364 64296 104364
rect 64495 100397 64613 104331
rect 64884 100364 64944 104364
rect 65144 100364 65216 104364
rect 65415 100397 65533 104331
rect 65804 100364 65864 104364
rect 66064 100364 66136 104364
rect 66335 100397 66453 104331
rect 66724 100364 66784 104364
rect 66984 100364 67056 104364
rect 67255 100397 67373 104331
rect 67644 100364 67704 104364
rect 67904 100364 67976 104364
rect 68175 100397 68293 104331
rect 68564 100364 68624 104364
rect 68824 100364 68896 104364
rect 69095 100397 69213 104331
rect 69484 100364 69544 104364
rect 80176 101334 80248 105334
rect 80447 101367 80565 105301
rect 80836 101334 80896 105334
rect 81096 101334 81168 105334
rect 81367 101367 81485 105301
rect 81756 101334 81816 105334
rect 82016 101334 82088 105334
rect 82287 101367 82405 105301
rect 82676 101334 82736 105334
rect 82936 101334 83008 105334
rect 83207 101367 83325 105301
rect 83596 101334 83656 105334
rect 83856 101334 83928 105334
rect 84127 101367 84245 105301
rect 84516 101334 84576 105334
rect 84776 101334 84848 105334
rect 85047 101367 85165 105301
rect 85436 101334 85496 105334
rect 85696 101334 85768 105334
rect 85967 101367 86085 105301
rect 86356 101334 86416 105334
rect 86616 101334 86688 105334
rect 86887 101367 87005 105301
rect 87276 101334 87336 105334
rect 87536 101334 87608 105334
rect 87807 101367 87925 105301
rect 88196 101334 88256 105334
rect 88456 101334 88528 105334
rect 88727 101367 88845 105301
rect 89116 101334 89176 105334
rect 89376 101334 89448 105334
rect 89647 101367 89765 105301
rect 90036 101334 90096 105334
rect 130062 105043 130112 105159
rect 130059 104959 130112 105043
rect 130232 104959 130360 105159
rect 130408 104959 130464 105159
rect 130584 104959 130712 105159
rect 130760 104959 130816 105159
rect 130936 104959 131064 105159
rect 131112 104959 131168 105159
rect 131288 104959 131416 105159
rect 131464 105043 131514 105159
rect 133925 105105 134925 105155
rect 131464 104959 131517 105043
rect 130067 104955 130101 104959
rect 131475 104955 131509 104959
rect 133925 104949 134925 105077
rect 133925 104793 134925 104921
rect 130000 104645 131000 104695
rect 132192 104645 133192 104695
rect 133925 104637 134925 104765
rect 122363 104026 122413 104626
rect 122513 104026 122563 104626
rect 122643 104026 122693 104626
rect 122793 104026 122921 104626
rect 122949 104026 123077 104626
rect 123105 104026 123161 104626
rect 123261 104026 123389 104626
rect 123417 104026 123545 104626
rect 123573 104026 123623 104626
rect 130000 104489 131000 104545
rect 132192 104489 133192 104545
rect 133925 104481 134925 104609
rect 131338 104405 131422 104408
rect 130000 104333 131000 104389
rect 131222 104355 131422 104405
rect 131770 104405 131854 104408
rect 131770 104400 131970 104405
rect 131766 104366 131970 104400
rect 131770 104355 131970 104366
rect 132192 104333 133192 104389
rect 133925 104325 134925 104453
rect 130000 104177 131000 104233
rect 131222 104179 131422 104307
rect 131770 104179 131970 104307
rect 132192 104177 133192 104233
rect 133925 104169 134925 104297
rect 130000 104021 131000 104077
rect 131222 104003 131422 104059
rect 131770 104003 131970 104059
rect 132192 104021 133192 104077
rect 133925 104013 134925 104141
rect 130000 103871 131000 103921
rect 130458 103868 130542 103871
rect 130790 103868 130874 103871
rect 131222 103827 131422 103955
rect 131770 103827 131970 103955
rect 132192 103871 133192 103921
rect 132318 103868 132402 103871
rect 132650 103868 132734 103871
rect 133925 103857 134925 103985
rect 99739 103696 99740 103720
rect 99820 103696 99821 103720
rect 100293 103696 100294 103720
rect 100374 103696 100375 103720
rect 100847 103696 100848 103720
rect 100928 103696 100929 103720
rect 101401 103696 101402 103720
rect 101482 103696 101483 103720
rect 101955 103696 101956 103720
rect 102036 103696 102037 103720
rect 102509 103696 102510 103720
rect 102590 103696 102591 103720
rect 103063 103696 103064 103720
rect 103144 103696 103145 103720
rect 103617 103696 103618 103720
rect 103698 103696 103699 103720
rect 104171 103696 104172 103720
rect 104252 103696 104253 103720
rect 104725 103696 104726 103720
rect 104806 103696 104807 103720
rect 105279 103696 105280 103720
rect 105360 103696 105361 103720
rect 105833 103696 105834 103720
rect 105914 103696 105915 103720
rect 106387 103696 106388 103720
rect 106468 103696 106469 103720
rect 106941 103696 106942 103720
rect 107022 103696 107023 103720
rect 107495 103696 107496 103720
rect 107576 103696 107577 103720
rect 108049 103696 108050 103720
rect 108130 103696 108131 103720
rect 108603 103696 108604 103720
rect 108684 103696 108685 103720
rect 109157 103696 109158 103720
rect 109238 103696 109239 103720
rect 109711 103696 109712 103720
rect 109792 103696 109793 103720
rect 110265 103696 110266 103720
rect 110346 103696 110347 103720
rect 99763 103672 99797 103684
rect 100317 103672 100351 103684
rect 100871 103672 100905 103684
rect 101425 103672 101459 103684
rect 101979 103672 102013 103684
rect 102533 103672 102567 103684
rect 103087 103672 103121 103684
rect 103641 103672 103675 103684
rect 104195 103672 104229 103684
rect 104749 103672 104783 103684
rect 105303 103672 105337 103684
rect 105857 103672 105891 103684
rect 106411 103672 106445 103684
rect 106965 103672 106999 103684
rect 107519 103672 107553 103684
rect 108073 103672 108107 103684
rect 108627 103672 108661 103684
rect 109181 103672 109215 103684
rect 109735 103672 109769 103684
rect 110289 103672 110323 103684
rect 125664 103634 125698 103668
rect 125733 103634 125767 103668
rect 125802 103634 125836 103668
rect 125871 103634 125905 103668
rect 125940 103634 125974 103668
rect 126009 103634 126043 103668
rect 126078 103634 126112 103668
rect 126147 103634 126181 103668
rect 126216 103634 126250 103668
rect 126285 103634 126319 103668
rect 126354 103634 126388 103668
rect 126423 103634 126457 103668
rect 126492 103634 126526 103668
rect 126561 103634 126595 103668
rect 126630 103634 126664 103668
rect 126699 103634 126733 103668
rect 126768 103634 126802 103668
rect 126837 103634 126871 103668
rect 126906 103634 126940 103668
rect 126975 103634 127009 103668
rect 127044 103634 127078 103668
rect 127113 103634 127147 103668
rect 127182 103634 127216 103668
rect 127251 103634 127285 103668
rect 127320 103634 127354 103668
rect 127389 103634 127423 103668
rect 127458 103634 127492 103668
rect 127527 103634 127561 103668
rect 127596 103634 127630 103668
rect 127665 103634 127699 103668
rect 127734 103635 127763 103668
rect 131222 103657 131422 103707
rect 131770 103657 131970 103707
rect 133925 103701 134925 103829
rect 127734 103634 127797 103635
rect 125664 103610 125688 103634
rect 133925 103545 134925 103673
rect 133925 103389 134925 103517
rect 133925 103233 134925 103361
rect 133925 103077 134925 103205
rect 133925 102927 134925 102977
rect 128376 102515 128400 102539
rect 128436 102515 128460 102539
rect 130751 102515 130775 102539
rect 130810 102515 130834 102539
rect 127858 102481 128306 102515
rect 128412 102491 128424 102515
rect 130786 102491 130799 102515
rect 130904 102481 131352 102515
rect 128414 102427 128448 102437
rect 128390 102416 128448 102427
rect 126030 102403 128448 102416
rect 130796 102416 130830 102437
rect 131423 102427 131457 102437
rect 131399 102416 131457 102427
rect 130796 102403 131457 102416
rect 126030 102395 128414 102403
rect 130796 102395 131423 102403
rect 133133 102402 133157 102426
rect 126030 102386 131613 102395
rect 133062 102386 133133 102392
rect 126030 102365 131583 102386
rect 133109 102378 133133 102386
rect 99739 101696 99740 101720
rect 99820 101696 99821 101720
rect 100293 101696 100294 101720
rect 100374 101696 100375 101720
rect 100847 101696 100848 101720
rect 100928 101696 100929 101720
rect 101401 101696 101402 101720
rect 101482 101696 101483 101720
rect 101955 101696 101956 101720
rect 102036 101696 102037 101720
rect 102509 101696 102510 101720
rect 102590 101696 102591 101720
rect 103063 101696 103064 101720
rect 103144 101696 103145 101720
rect 103617 101696 103618 101720
rect 103698 101696 103699 101720
rect 104171 101696 104172 101720
rect 104252 101696 104253 101720
rect 104725 101696 104726 101720
rect 104806 101696 104807 101720
rect 105279 101696 105280 101720
rect 105360 101696 105361 101720
rect 105833 101696 105834 101720
rect 105914 101696 105915 101720
rect 106387 101696 106388 101720
rect 106468 101696 106469 101720
rect 106941 101696 106942 101720
rect 107022 101696 107023 101720
rect 107495 101696 107496 101720
rect 107576 101696 107577 101720
rect 108049 101696 108050 101720
rect 108130 101696 108131 101720
rect 108603 101696 108604 101720
rect 108684 101696 108685 101720
rect 109157 101696 109158 101720
rect 109238 101696 109239 101720
rect 109711 101696 109712 101720
rect 109792 101696 109793 101720
rect 110265 101696 110266 101720
rect 110346 101696 110347 101720
rect 99763 101672 99797 101684
rect 100317 101672 100351 101684
rect 100871 101672 100905 101684
rect 101425 101672 101459 101684
rect 101979 101672 102013 101684
rect 102533 101672 102567 101684
rect 103087 101672 103121 101684
rect 103641 101672 103675 101684
rect 104195 101672 104229 101684
rect 104749 101672 104783 101684
rect 105303 101672 105337 101684
rect 105857 101672 105891 101684
rect 106411 101672 106445 101684
rect 106965 101672 106999 101684
rect 107519 101672 107553 101684
rect 108073 101672 108107 101684
rect 108627 101672 108661 101684
rect 109181 101672 109215 101684
rect 109735 101672 109769 101684
rect 110289 101672 110323 101684
rect 121250 101546 121300 102146
rect 121420 101546 121476 102146
rect 121596 101546 121646 102146
rect 119951 101460 119975 101484
rect 120012 101474 120036 101484
rect 120012 101470 120046 101474
rect 120083 101470 120117 101474
rect 120154 101470 120188 101474
rect 119990 101460 120212 101470
rect 119988 101456 119999 101460
rect 120012 101456 120046 101460
rect 120083 101456 120117 101460
rect 120154 101456 120188 101460
rect 119988 101436 120212 101456
rect 120012 101416 120036 101436
rect 121735 101324 121785 102324
rect 121885 101324 121935 102324
rect 122044 101324 122094 102324
rect 122194 101324 122244 102324
rect 122374 101864 122554 102064
rect 122719 102049 122779 102064
rect 122805 102049 122865 102064
rect 124379 102049 124439 102064
rect 124465 102049 124525 102064
rect 122734 101879 122764 102049
rect 122820 101879 122850 102049
rect 124394 101879 124424 102049
rect 124480 101879 124510 102049
rect 122723 101876 122775 101879
rect 122809 101876 122861 101879
rect 124383 101876 124435 101879
rect 124469 101876 124521 101879
rect 122719 101864 122779 101876
rect 122805 101864 122865 101876
rect 124379 101864 124439 101876
rect 124465 101864 124525 101876
rect 124690 101864 124870 102064
rect 122374 101604 122554 101804
rect 122719 101789 122779 101804
rect 122805 101789 122865 101804
rect 124379 101789 124439 101804
rect 124465 101789 124525 101804
rect 122734 101619 122764 101789
rect 122820 101619 122850 101789
rect 124394 101619 124424 101789
rect 124480 101619 124510 101789
rect 122723 101616 122775 101619
rect 122809 101616 122861 101619
rect 124383 101616 124435 101619
rect 124469 101616 124521 101619
rect 122719 101604 122779 101616
rect 122805 101604 122865 101616
rect 124379 101604 124439 101616
rect 124465 101604 124525 101616
rect 124690 101604 124870 101804
rect 122374 101344 122554 101544
rect 122719 101529 122779 101544
rect 122805 101529 122865 101544
rect 124379 101529 124439 101544
rect 124465 101529 124525 101544
rect 122734 101524 122764 101529
rect 122820 101524 122850 101529
rect 124394 101524 124424 101529
rect 124480 101524 124510 101529
rect 124690 101344 124870 101544
rect 125000 101324 125050 102324
rect 125150 101324 125200 102324
rect 125309 101324 125359 102324
rect 125459 101324 125509 102324
rect 126787 102302 132608 102338
rect 126787 102290 126823 102302
rect 126873 102290 126907 102302
rect 126942 102290 126976 102302
rect 127011 102290 127045 102302
rect 127080 102290 127114 102302
rect 127149 102290 127183 102302
rect 127218 102290 127252 102302
rect 127287 102290 127321 102302
rect 127356 102290 127390 102302
rect 127425 102290 127459 102302
rect 127494 102290 127528 102302
rect 127563 102290 127597 102302
rect 127632 102290 127666 102302
rect 127701 102290 127735 102302
rect 127770 102290 127804 102302
rect 127839 102290 127873 102302
rect 127908 102290 127942 102302
rect 127977 102290 128011 102302
rect 128046 102290 128080 102302
rect 128115 102290 128149 102302
rect 128184 102290 128218 102302
rect 128253 102290 128287 102302
rect 128322 102290 128356 102302
rect 128391 102290 128425 102302
rect 128460 102290 128494 102302
rect 128529 102290 128563 102302
rect 128598 102290 128632 102302
rect 128667 102290 128701 102302
rect 128736 102290 128770 102302
rect 128805 102290 128839 102302
rect 128874 102290 128908 102302
rect 128943 102290 128977 102302
rect 129012 102290 129046 102302
rect 129081 102290 129115 102302
rect 129150 102290 129184 102302
rect 129219 102290 129253 102302
rect 129288 102290 129322 102302
rect 129357 102290 129391 102302
rect 129426 102290 129460 102302
rect 129495 102290 129529 102302
rect 129564 102290 129598 102302
rect 129633 102290 129667 102302
rect 129702 102290 129736 102302
rect 129771 102290 129805 102302
rect 129840 102290 129874 102302
rect 129909 102290 129943 102302
rect 129978 102290 130012 102302
rect 130047 102290 130081 102302
rect 130116 102290 130150 102302
rect 130185 102290 130219 102302
rect 130254 102290 130288 102302
rect 130323 102290 130357 102302
rect 130392 102290 130426 102302
rect 130461 102290 130495 102302
rect 130530 102290 130564 102302
rect 130599 102290 130633 102302
rect 130668 102290 130702 102302
rect 130737 102290 130771 102302
rect 130806 102290 130840 102302
rect 130875 102290 130909 102302
rect 130944 102290 130978 102302
rect 131013 102290 131047 102302
rect 131082 102290 131116 102302
rect 131151 102290 131185 102302
rect 131220 102290 131254 102302
rect 131289 102290 131323 102302
rect 131358 102290 131392 102302
rect 131426 102290 131460 102302
rect 131494 102290 131528 102302
rect 131562 102290 131596 102302
rect 131630 102290 131664 102302
rect 131698 102290 131732 102302
rect 131766 102290 131800 102302
rect 131834 102290 131868 102302
rect 131902 102290 131936 102302
rect 131970 102290 132004 102302
rect 132038 102290 132072 102302
rect 132106 102290 132140 102302
rect 132174 102290 132208 102302
rect 132242 102290 132276 102302
rect 132310 102290 132344 102302
rect 132378 102290 132412 102302
rect 132446 102290 132480 102302
rect 132514 102290 132548 102302
rect 132572 102290 132608 102302
rect 126787 102254 126839 102290
rect 125598 101546 125648 102146
rect 125768 101546 125824 102146
rect 125944 101546 125994 102146
rect 126823 101599 126839 102254
rect 126803 101596 126839 101599
rect 126849 101596 126885 102290
rect 126907 102254 126942 102290
rect 126976 102254 127011 102290
rect 127045 102254 127080 102290
rect 127114 102254 127149 102290
rect 127183 102254 127218 102290
rect 127252 102254 127287 102290
rect 127321 102254 127356 102290
rect 127390 102254 127425 102290
rect 127459 102254 127494 102290
rect 127528 102254 127563 102290
rect 127597 102254 127632 102290
rect 127666 102254 127701 102290
rect 127735 102254 127770 102290
rect 127804 102254 127839 102290
rect 127873 102254 127908 102290
rect 127942 102254 127977 102290
rect 128011 102254 128046 102290
rect 128080 102254 128115 102290
rect 128149 102254 128184 102290
rect 128218 102254 128253 102290
rect 128287 102254 128322 102290
rect 128356 102254 128391 102290
rect 128425 102254 128460 102290
rect 128494 102254 128529 102290
rect 128563 102254 128598 102290
rect 128632 102254 128667 102290
rect 128701 102254 128736 102290
rect 128770 102254 128805 102290
rect 128839 102254 128874 102290
rect 128908 102254 128943 102290
rect 128977 102254 129012 102290
rect 129046 102254 129081 102290
rect 129115 102254 129150 102290
rect 129184 102254 129219 102290
rect 129253 102254 129288 102290
rect 129322 102254 129357 102290
rect 129391 102254 129426 102290
rect 129460 102254 129495 102290
rect 129529 102254 129564 102290
rect 129598 102254 129633 102290
rect 129667 102254 129702 102290
rect 129736 102254 129771 102290
rect 129805 102254 129840 102290
rect 129874 102254 129909 102290
rect 129943 102254 129978 102290
rect 130012 102254 130047 102290
rect 130081 102254 130116 102290
rect 130150 102254 130185 102290
rect 130219 102254 130254 102290
rect 130288 102254 130323 102290
rect 130357 102254 130392 102290
rect 130426 102254 130461 102290
rect 130495 102254 130530 102290
rect 130564 102254 130599 102290
rect 130633 102254 130668 102290
rect 130702 102254 130737 102290
rect 130771 102254 130806 102290
rect 130840 102254 130875 102290
rect 130909 102254 130944 102290
rect 130978 102254 131013 102290
rect 131047 102254 131082 102290
rect 131116 102254 131151 102290
rect 131185 102254 131220 102290
rect 131254 102254 131289 102290
rect 131323 102254 131358 102290
rect 131392 102254 131426 102290
rect 131460 102254 131494 102290
rect 131528 102254 131562 102290
rect 131596 102254 131630 102290
rect 131664 102254 131698 102290
rect 131732 102254 131766 102290
rect 131800 102254 131834 102290
rect 131868 102254 131902 102290
rect 131936 102254 131970 102290
rect 132004 102254 132038 102290
rect 132072 102254 132106 102290
rect 132140 102254 132174 102290
rect 132208 102254 132242 102290
rect 132276 102254 132310 102290
rect 132344 102254 132378 102290
rect 132412 102254 132446 102290
rect 132480 102254 132514 102290
rect 132548 102254 132608 102290
rect 126803 101560 126885 101596
rect 126983 101582 127033 102182
rect 127153 101582 127209 102182
rect 127329 101582 127379 102182
rect 127445 101582 127495 102182
rect 127615 101582 127671 102182
rect 127791 101582 127919 102182
rect 127967 101582 128095 102182
rect 128143 101582 128271 102182
rect 128319 101582 128369 102182
rect 128435 101582 128485 102182
rect 128605 101582 128733 102182
rect 128781 101582 128837 102182
rect 128957 101582 129085 102182
rect 129133 101582 129183 102182
rect 129249 101582 129299 102182
rect 129419 101582 129547 102182
rect 129595 101582 129723 102182
rect 129771 101582 129899 102182
rect 129947 101582 130075 102182
rect 130123 101582 130251 102182
rect 130299 101582 130355 102182
rect 130475 101582 130603 102182
rect 130651 101582 130779 102182
rect 130827 101582 130955 102182
rect 131003 101582 131131 102182
rect 131179 101582 131307 102182
rect 131355 101582 131411 102182
rect 131531 101582 131659 102182
rect 131707 101582 131763 102182
rect 131883 101582 132011 102182
rect 132059 101582 132115 102182
rect 132235 101582 132363 102182
rect 132411 101582 132461 102182
rect 133886 101872 134066 102072
rect 134122 101872 134302 102072
rect 133886 101737 134066 101774
rect 134573 101472 134623 102072
rect 134743 101472 134799 102072
rect 134919 101472 134975 102072
rect 135095 101472 135145 102072
rect 122374 101030 122554 101230
rect 124690 101030 124870 101230
rect 120738 100254 120788 100854
rect 120888 100254 120944 100854
rect 121044 100254 121094 100854
rect 121778 100770 121958 100970
rect 122014 100770 122194 100970
rect 122374 100770 122554 100970
rect 122719 100955 122779 100970
rect 122805 100955 122865 100970
rect 124379 100955 124439 100970
rect 124465 100955 124525 100970
rect 122734 100785 122764 100955
rect 122820 100785 122850 100955
rect 122975 100836 123063 100872
rect 122975 100832 123011 100836
rect 123027 100832 123063 100836
rect 123011 100798 123063 100832
rect 122723 100782 122775 100785
rect 122809 100782 122861 100785
rect 122719 100770 122779 100782
rect 122805 100770 122865 100782
rect 122975 100764 123011 100798
rect 123027 100764 123063 100798
rect 123011 100730 123063 100764
rect 121778 100510 121958 100710
rect 122014 100510 122194 100710
rect 122374 100510 122554 100710
rect 122719 100695 122779 100710
rect 122805 100695 122865 100710
rect 122975 100696 123011 100730
rect 123027 100696 123063 100730
rect 122734 100525 122764 100695
rect 122820 100525 122850 100695
rect 123011 100662 123063 100696
rect 122975 100628 123011 100662
rect 123027 100628 123063 100662
rect 123011 100594 123063 100628
rect 122975 100560 123011 100594
rect 123027 100560 123063 100594
rect 123011 100526 123063 100560
rect 122723 100522 122775 100525
rect 122809 100522 122861 100525
rect 122719 100510 122779 100522
rect 122805 100510 122865 100522
rect 122975 100494 123011 100526
rect 123027 100520 123063 100526
rect 122374 100250 122554 100450
rect 122719 100435 122779 100450
rect 122805 100435 122865 100450
rect 122734 100396 122764 100435
rect 122820 100396 122850 100435
rect 122977 100256 123011 100494
rect 123015 100484 123063 100520
rect 124179 100836 124269 100872
rect 124179 100520 124215 100836
rect 124233 100520 124269 100836
rect 124394 100785 124424 100955
rect 124480 100785 124510 100955
rect 124383 100782 124435 100785
rect 124469 100782 124521 100785
rect 124379 100770 124439 100782
rect 124465 100770 124525 100782
rect 124690 100770 124870 100970
rect 125050 100770 125230 100970
rect 125286 100770 125466 100970
rect 124379 100695 124439 100710
rect 124465 100695 124525 100710
rect 124394 100525 124424 100695
rect 124480 100525 124510 100695
rect 124383 100522 124435 100525
rect 124469 100522 124521 100525
rect 124179 100484 124269 100520
rect 124379 100510 124439 100522
rect 124465 100510 124525 100522
rect 124690 100510 124870 100710
rect 125050 100510 125230 100710
rect 125286 100510 125466 100710
rect 123015 100256 123051 100484
rect 124235 100256 124267 100484
rect 124379 100435 124439 100450
rect 124465 100435 124525 100450
rect 124394 100396 124424 100435
rect 124480 100396 124510 100435
rect 122975 100220 123051 100256
rect 124690 100250 124870 100450
rect 126150 100254 126200 100854
rect 126300 100254 126356 100854
rect 126456 100254 126506 100854
rect 127003 100268 127053 101268
rect 127153 100268 127209 101268
rect 127309 100268 127359 101268
rect 127445 100268 127495 101268
rect 127595 100268 127651 101268
rect 127751 100268 127807 101268
rect 127907 100268 127963 101268
rect 128063 100268 128113 101268
rect 128179 100268 128229 101268
rect 128329 100268 128457 101268
rect 128485 100268 128613 101268
rect 128641 100268 128769 101268
rect 128797 100268 128925 101268
rect 128953 100268 129081 101268
rect 129109 100268 129165 101268
rect 129265 100268 129393 101268
rect 129421 100268 129549 101268
rect 129577 100268 129705 101268
rect 129733 100268 129861 101268
rect 129889 100268 130017 101268
rect 130045 100268 130101 101268
rect 130221 100268 130349 101268
rect 130397 100268 130525 101268
rect 130573 100268 130701 101268
rect 130749 100268 130877 101268
rect 130925 100268 131053 101268
rect 131101 100268 131229 101268
rect 131277 100268 131405 101268
rect 131453 100268 131503 101268
rect 131569 100268 131619 101268
rect 131719 100268 131847 101268
rect 131875 100268 132003 101268
rect 132031 100268 132159 101268
rect 132187 100268 132243 101268
rect 132343 100268 132471 101268
rect 132499 100268 132627 101268
rect 132655 100268 132783 101268
rect 132811 100268 132861 101268
rect 133452 100709 133505 100859
rect 133455 100612 133505 100709
rect 133452 100390 133505 100612
rect 133455 100259 133505 100390
rect 133625 100259 133681 100859
rect 133801 100259 133851 100859
rect 134227 100264 134277 100864
rect 134397 100264 134447 100864
rect 1823 99308 1824 99332
rect 1904 99308 1905 99332
rect 2377 99308 2378 99332
rect 2458 99308 2459 99332
rect 2931 99308 2932 99332
rect 3012 99308 3013 99332
rect 3485 99308 3486 99332
rect 3566 99308 3567 99332
rect 4039 99308 4040 99332
rect 4120 99308 4121 99332
rect 4593 99308 4594 99332
rect 4674 99308 4675 99332
rect 5147 99308 5148 99332
rect 5228 99308 5229 99332
rect 5701 99308 5702 99332
rect 5782 99308 5783 99332
rect 6255 99308 6256 99332
rect 6336 99308 6337 99332
rect 6809 99308 6810 99332
rect 6890 99308 6891 99332
rect 7363 99308 7364 99332
rect 7444 99308 7445 99332
rect 7917 99308 7918 99332
rect 7998 99308 7999 99332
rect 8471 99308 8472 99332
rect 8552 99308 8553 99332
rect 9025 99308 9026 99332
rect 9106 99308 9107 99332
rect 9579 99308 9580 99332
rect 9660 99308 9661 99332
rect 10133 99308 10134 99332
rect 10214 99308 10215 99332
rect 10687 99308 10688 99332
rect 10768 99308 10769 99332
rect 11241 99308 11242 99332
rect 11322 99308 11323 99332
rect 11795 99308 11796 99332
rect 11876 99308 11877 99332
rect 12349 99308 12350 99332
rect 12430 99308 12431 99332
rect 1847 99284 1881 99296
rect 2401 99284 2435 99296
rect 2955 99284 2989 99296
rect 3509 99284 3543 99296
rect 4063 99284 4097 99296
rect 4617 99284 4651 99296
rect 5171 99284 5205 99296
rect 5725 99284 5759 99296
rect 6279 99284 6313 99296
rect 6833 99284 6867 99296
rect 7387 99284 7421 99296
rect 7941 99284 7975 99296
rect 8495 99284 8529 99296
rect 9049 99284 9083 99296
rect 9603 99284 9637 99296
rect 10157 99284 10191 99296
rect 10711 99284 10745 99296
rect 11265 99284 11299 99296
rect 11819 99284 11853 99296
rect 12373 99284 12407 99296
rect 20904 98024 20954 99424
rect 21054 98024 21182 99424
rect 21210 98024 21338 99424
rect 21366 98024 21494 99424
rect 21522 98024 21650 99424
rect 21678 98024 21806 99424
rect 21834 98024 21962 99424
rect 21990 98024 22118 99424
rect 22146 98024 22274 99424
rect 22302 98024 22430 99424
rect 22458 98024 22586 99424
rect 22614 98024 22742 99424
rect 22770 98024 22898 99424
rect 22926 98024 23054 99424
rect 23082 98024 23210 99424
rect 23238 98024 23366 99424
rect 23394 98024 23522 99424
rect 23550 98024 23678 99424
rect 23706 98024 23834 99424
rect 23862 98024 23990 99424
rect 24018 98024 24146 99424
rect 24174 98024 24302 99424
rect 24330 98024 24458 99424
rect 24486 98024 24614 99424
rect 24642 98024 24770 99424
rect 24798 98024 24926 99424
rect 24954 98024 25082 99424
rect 25110 98024 25238 99424
rect 25266 98024 25394 99424
rect 25422 98024 25550 99424
rect 25578 98024 25706 99424
rect 25734 98024 25862 99424
rect 25890 98024 26018 99424
rect 26046 98024 26174 99424
rect 26202 98024 26330 99424
rect 26358 98024 26486 99424
rect 26514 98024 26642 99424
rect 26670 98024 26798 99424
rect 26826 98024 26954 99424
rect 26982 98024 27110 99424
rect 27138 98024 27266 99424
rect 27294 98024 27422 99424
rect 27450 98024 27578 99424
rect 27606 98024 27734 99424
rect 27762 98024 27890 99424
rect 27918 98024 28046 99424
rect 28074 98024 28202 99424
rect 28230 98024 28358 99424
rect 28386 98024 28514 99424
rect 28542 98024 28670 99424
rect 28698 98024 28748 99424
rect 30619 98580 30669 99980
rect 30769 98580 30897 99980
rect 30925 98580 31053 99980
rect 31081 98580 31209 99980
rect 31237 98580 31365 99980
rect 31393 98580 31521 99980
rect 31549 98580 31677 99980
rect 31705 98580 31833 99980
rect 31861 98580 31989 99980
rect 32017 98580 32145 99980
rect 32173 98580 32301 99980
rect 32329 98580 32457 99980
rect 32485 98580 32613 99980
rect 32641 98580 32769 99980
rect 32797 98580 32925 99980
rect 32953 98580 33003 99980
rect 40797 98532 40798 98556
rect 40878 98532 40879 98556
rect 41351 98532 41352 98556
rect 41432 98532 41433 98556
rect 41905 98532 41906 98556
rect 41986 98532 41987 98556
rect 42459 98532 42460 98556
rect 42540 98532 42541 98556
rect 43013 98532 43014 98556
rect 43094 98532 43095 98556
rect 43567 98532 43568 98556
rect 43648 98532 43649 98556
rect 44121 98532 44122 98556
rect 44202 98532 44203 98556
rect 44675 98532 44676 98556
rect 44756 98532 44757 98556
rect 45229 98532 45230 98556
rect 45310 98532 45311 98556
rect 45783 98532 45784 98556
rect 45864 98532 45865 98556
rect 46337 98532 46338 98556
rect 46418 98532 46419 98556
rect 46891 98532 46892 98556
rect 46972 98532 46973 98556
rect 47445 98532 47446 98556
rect 47526 98532 47527 98556
rect 47999 98532 48000 98556
rect 48080 98532 48081 98556
rect 48553 98532 48554 98556
rect 48634 98532 48635 98556
rect 49107 98532 49108 98556
rect 49188 98532 49189 98556
rect 49661 98532 49662 98556
rect 49742 98532 49743 98556
rect 50215 98532 50216 98556
rect 50296 98532 50297 98556
rect 50769 98532 50770 98556
rect 50850 98532 50851 98556
rect 51323 98532 51324 98556
rect 51404 98532 51405 98556
rect 40821 98508 40855 98520
rect 41375 98508 41409 98520
rect 41929 98508 41963 98520
rect 42483 98508 42517 98520
rect 43037 98508 43071 98520
rect 43591 98508 43625 98520
rect 44145 98508 44179 98520
rect 44699 98508 44733 98520
rect 45253 98508 45287 98520
rect 45807 98508 45841 98520
rect 46361 98508 46395 98520
rect 46915 98508 46949 98520
rect 47469 98508 47503 98520
rect 48023 98508 48057 98520
rect 48577 98508 48611 98520
rect 49131 98508 49165 98520
rect 49685 98508 49719 98520
rect 50239 98508 50273 98520
rect 50793 98508 50827 98520
rect 51347 98508 51381 98520
rect 1823 97308 1824 97332
rect 1904 97308 1905 97332
rect 2377 97308 2378 97332
rect 2458 97308 2459 97332
rect 2931 97308 2932 97332
rect 3012 97308 3013 97332
rect 3485 97308 3486 97332
rect 3566 97308 3567 97332
rect 4039 97308 4040 97332
rect 4120 97308 4121 97332
rect 4593 97308 4594 97332
rect 4674 97308 4675 97332
rect 5147 97308 5148 97332
rect 5228 97308 5229 97332
rect 5701 97308 5702 97332
rect 5782 97308 5783 97332
rect 6255 97308 6256 97332
rect 6336 97308 6337 97332
rect 6809 97308 6810 97332
rect 6890 97308 6891 97332
rect 7363 97308 7364 97332
rect 7444 97308 7445 97332
rect 7917 97308 7918 97332
rect 7998 97308 7999 97332
rect 8471 97308 8472 97332
rect 8552 97308 8553 97332
rect 9025 97308 9026 97332
rect 9106 97308 9107 97332
rect 9579 97308 9580 97332
rect 9660 97308 9661 97332
rect 10133 97308 10134 97332
rect 10214 97308 10215 97332
rect 10687 97308 10688 97332
rect 10768 97308 10769 97332
rect 11241 97308 11242 97332
rect 11322 97308 11323 97332
rect 11795 97308 11796 97332
rect 11876 97308 11877 97332
rect 12349 97308 12350 97332
rect 12430 97308 12431 97332
rect 1847 97284 1881 97296
rect 2401 97284 2435 97296
rect 2955 97284 2989 97296
rect 3509 97284 3543 97296
rect 4063 97284 4097 97296
rect 4617 97284 4651 97296
rect 5171 97284 5205 97296
rect 5725 97284 5759 97296
rect 6279 97284 6313 97296
rect 6833 97284 6867 97296
rect 7387 97284 7421 97296
rect 7941 97284 7975 97296
rect 8495 97284 8529 97296
rect 9049 97284 9083 97296
rect 9603 97284 9637 97296
rect 10157 97284 10191 97296
rect 10711 97284 10745 97296
rect 11265 97284 11299 97296
rect 11819 97284 11853 97296
rect 12373 97284 12407 97296
rect 31199 96493 31249 97493
rect 32049 96493 32099 97493
rect 32351 96493 32401 97493
rect 33201 96493 33251 97493
rect 57744 96888 57794 98288
rect 57894 96888 58022 98288
rect 58050 96888 58178 98288
rect 58206 96888 58334 98288
rect 58362 96888 58490 98288
rect 58518 96888 58646 98288
rect 58674 96888 58802 98288
rect 58830 96888 58958 98288
rect 58986 96888 59114 98288
rect 59142 96888 59270 98288
rect 59298 96888 59426 98288
rect 59454 96888 59582 98288
rect 59610 96888 59738 98288
rect 59766 96888 59894 98288
rect 59922 96888 60050 98288
rect 60078 96888 60206 98288
rect 60234 96888 60362 98288
rect 60390 96888 60518 98288
rect 60546 96888 60674 98288
rect 60702 96888 60830 98288
rect 60858 96888 60986 98288
rect 61014 96888 61142 98288
rect 61170 96888 61298 98288
rect 61326 96888 61454 98288
rect 61482 96888 61610 98288
rect 61638 96888 61766 98288
rect 61794 96888 61922 98288
rect 61950 96888 62078 98288
rect 62106 96888 62234 98288
rect 62262 96888 62390 98288
rect 62418 96888 62546 98288
rect 62574 96888 62702 98288
rect 62730 96888 62858 98288
rect 62886 96888 63014 98288
rect 63042 96888 63170 98288
rect 63198 96888 63326 98288
rect 63354 96888 63482 98288
rect 63510 96888 63638 98288
rect 63666 96888 63794 98288
rect 63822 96888 63950 98288
rect 63978 96888 64106 98288
rect 64134 96888 64262 98288
rect 64290 96888 64418 98288
rect 64446 96888 64574 98288
rect 64602 96888 64730 98288
rect 64758 96888 64886 98288
rect 64914 96888 65042 98288
rect 65070 96888 65198 98288
rect 65226 96888 65354 98288
rect 65382 96888 65510 98288
rect 65538 96888 65588 98288
rect 67459 97444 67509 98844
rect 67609 97444 67737 98844
rect 67765 97444 67893 98844
rect 67921 97444 68049 98844
rect 68077 97444 68205 98844
rect 68233 97444 68361 98844
rect 68389 97444 68517 98844
rect 68545 97444 68673 98844
rect 68701 97444 68829 98844
rect 68857 97444 68985 98844
rect 69013 97444 69141 98844
rect 69169 97444 69297 98844
rect 69325 97444 69453 98844
rect 69481 97444 69609 98844
rect 69637 97444 69765 98844
rect 69793 97444 69843 98844
rect 78296 97858 78346 99258
rect 78446 97858 78574 99258
rect 78602 97858 78730 99258
rect 78758 97858 78886 99258
rect 78914 97858 79042 99258
rect 79070 97858 79198 99258
rect 79226 97858 79354 99258
rect 79382 97858 79510 99258
rect 79538 97858 79666 99258
rect 79694 97858 79822 99258
rect 79850 97858 79978 99258
rect 80006 97858 80134 99258
rect 80162 97858 80290 99258
rect 80318 97858 80446 99258
rect 80474 97858 80602 99258
rect 80630 97858 80758 99258
rect 80786 97858 80914 99258
rect 80942 97858 81070 99258
rect 81098 97858 81226 99258
rect 81254 97858 81382 99258
rect 81410 97858 81538 99258
rect 81566 97858 81694 99258
rect 81722 97858 81850 99258
rect 81878 97858 82006 99258
rect 82034 97858 82162 99258
rect 82190 97858 82318 99258
rect 82346 97858 82474 99258
rect 82502 97858 82630 99258
rect 82658 97858 82786 99258
rect 82814 97858 82942 99258
rect 82970 97858 83098 99258
rect 83126 97858 83254 99258
rect 83282 97858 83410 99258
rect 83438 97858 83566 99258
rect 83594 97858 83722 99258
rect 83750 97858 83878 99258
rect 83906 97858 84034 99258
rect 84062 97858 84190 99258
rect 84218 97858 84346 99258
rect 84374 97858 84502 99258
rect 84530 97858 84658 99258
rect 84686 97858 84814 99258
rect 84842 97858 84970 99258
rect 84998 97858 85126 99258
rect 85154 97858 85282 99258
rect 85310 97858 85438 99258
rect 85466 97858 85594 99258
rect 85622 97858 85750 99258
rect 85778 97858 85906 99258
rect 85934 97858 86062 99258
rect 86090 97858 86140 99258
rect 88011 98414 88061 99814
rect 88161 98414 88289 99814
rect 88317 98414 88445 99814
rect 88473 98414 88601 99814
rect 88629 98414 88757 99814
rect 88785 98414 88913 99814
rect 88941 98414 89069 99814
rect 89097 98414 89225 99814
rect 89253 98414 89381 99814
rect 89409 98414 89537 99814
rect 89565 98414 89693 99814
rect 89721 98414 89849 99814
rect 89877 98414 90005 99814
rect 90033 98414 90161 99814
rect 90189 98414 90317 99814
rect 90345 98414 90395 99814
rect 99739 99696 99740 99720
rect 99820 99696 99821 99720
rect 100293 99696 100294 99720
rect 100374 99696 100375 99720
rect 100847 99696 100848 99720
rect 100928 99696 100929 99720
rect 101401 99696 101402 99720
rect 101482 99696 101483 99720
rect 101955 99696 101956 99720
rect 102036 99696 102037 99720
rect 102509 99696 102510 99720
rect 102590 99696 102591 99720
rect 103063 99696 103064 99720
rect 103144 99696 103145 99720
rect 103617 99696 103618 99720
rect 103698 99696 103699 99720
rect 104171 99696 104172 99720
rect 104252 99696 104253 99720
rect 104725 99696 104726 99720
rect 104806 99696 104807 99720
rect 105279 99696 105280 99720
rect 105360 99696 105361 99720
rect 105833 99696 105834 99720
rect 105914 99696 105915 99720
rect 106387 99696 106388 99720
rect 106468 99696 106469 99720
rect 106941 99696 106942 99720
rect 107022 99696 107023 99720
rect 107495 99696 107496 99720
rect 107576 99696 107577 99720
rect 108049 99696 108050 99720
rect 108130 99696 108131 99720
rect 108603 99696 108604 99720
rect 108684 99696 108685 99720
rect 109157 99696 109158 99720
rect 109238 99696 109239 99720
rect 109711 99696 109712 99720
rect 109792 99696 109793 99720
rect 110265 99696 110266 99720
rect 110346 99696 110347 99720
rect 99763 99672 99797 99684
rect 100317 99672 100351 99684
rect 100871 99672 100905 99684
rect 101425 99672 101459 99684
rect 101979 99672 102013 99684
rect 102533 99672 102567 99684
rect 103087 99672 103121 99684
rect 103641 99672 103675 99684
rect 104195 99672 104229 99684
rect 104749 99672 104783 99684
rect 105303 99672 105337 99684
rect 105857 99672 105891 99684
rect 106411 99672 106445 99684
rect 106965 99672 106999 99684
rect 107519 99672 107553 99684
rect 108073 99672 108107 99684
rect 108627 99672 108661 99684
rect 109181 99672 109215 99684
rect 109735 99672 109769 99684
rect 110289 99672 110323 99684
rect 119455 99282 119463 99507
rect 119532 98425 119582 99025
rect 119682 98425 119732 99025
rect 120588 98787 120638 99387
rect 120738 98787 120794 99387
rect 120894 98787 120944 99387
rect 121116 98721 121166 99721
rect 121266 98721 121322 99721
rect 121422 98721 121472 99721
rect 121538 98721 121588 99721
rect 121688 98721 121816 99721
rect 121844 98721 121972 99721
rect 122000 98721 122128 99721
rect 122156 98721 122212 99721
rect 122312 98721 122440 99721
rect 122468 98721 122596 99721
rect 122624 98721 122752 99721
rect 122780 98721 122830 99721
rect 122982 98721 123032 99721
rect 123132 98721 123260 99721
rect 123288 98721 123416 99721
rect 123444 98721 123572 99721
rect 123600 98721 123728 99721
rect 123756 98721 123884 99721
rect 123912 98721 124040 99721
rect 124068 98721 124196 99721
rect 124224 98721 124274 99721
rect 124426 98771 124476 99771
rect 124576 98771 124704 99771
rect 124732 98771 124860 99771
rect 124888 98771 125016 99771
rect 125044 98771 125172 99771
rect 125200 98771 125328 99771
rect 125356 98771 125484 99771
rect 125512 98771 125640 99771
rect 125668 98771 125718 99771
rect 125870 98721 125920 99721
rect 126020 98721 126148 99721
rect 126176 98721 126304 99721
rect 126332 98721 126460 99721
rect 126488 98721 126616 99721
rect 126644 98721 126772 99721
rect 126800 98721 126928 99721
rect 126956 98721 127084 99721
rect 127112 98721 127168 99721
rect 127268 98721 127318 99721
rect 127470 99121 127520 99721
rect 127904 99121 127954 99721
rect 129147 99236 129197 99836
rect 129297 99236 129425 99836
rect 129453 99236 129581 99836
rect 129609 99236 129659 99836
rect 129739 99236 129789 99836
rect 129889 99236 130017 99836
rect 130045 99236 130101 99836
rect 130201 99236 130329 99836
rect 130357 99236 130407 99836
rect 130487 99236 130537 99836
rect 130637 99236 130693 99836
rect 130793 99236 130843 99836
rect 129772 98456 129808 99056
rect 130132 98456 130188 99056
rect 130322 98456 130372 99056
rect 126035 98342 126101 98358
rect 126197 98342 126263 98358
rect 128605 98288 128680 98298
rect 128900 98288 128975 98298
rect 99739 97696 99740 97720
rect 99820 97696 99821 97720
rect 100293 97696 100294 97720
rect 100374 97696 100375 97720
rect 100847 97696 100848 97720
rect 100928 97696 100929 97720
rect 101401 97696 101402 97720
rect 101482 97696 101483 97720
rect 101955 97696 101956 97720
rect 102036 97696 102037 97720
rect 102509 97696 102510 97720
rect 102590 97696 102591 97720
rect 103063 97696 103064 97720
rect 103144 97696 103145 97720
rect 103617 97696 103618 97720
rect 103698 97696 103699 97720
rect 104171 97696 104172 97720
rect 104252 97696 104253 97720
rect 104725 97696 104726 97720
rect 104806 97696 104807 97720
rect 105279 97696 105280 97720
rect 105360 97696 105361 97720
rect 105833 97696 105834 97720
rect 105914 97696 105915 97720
rect 106387 97696 106388 97720
rect 106468 97696 106469 97720
rect 106941 97696 106942 97720
rect 107022 97696 107023 97720
rect 107495 97696 107496 97720
rect 107576 97696 107577 97720
rect 108049 97696 108050 97720
rect 108130 97696 108131 97720
rect 108603 97696 108604 97720
rect 108684 97696 108685 97720
rect 109157 97696 109158 97720
rect 109238 97696 109239 97720
rect 109711 97696 109712 97720
rect 109792 97696 109793 97720
rect 110265 97696 110266 97720
rect 110346 97696 110347 97720
rect 99763 97672 99797 97684
rect 100317 97672 100351 97684
rect 100871 97672 100905 97684
rect 101425 97672 101459 97684
rect 101979 97672 102013 97684
rect 102533 97672 102567 97684
rect 103087 97672 103121 97684
rect 103641 97672 103675 97684
rect 104195 97672 104229 97684
rect 104749 97672 104783 97684
rect 105303 97672 105337 97684
rect 105857 97672 105891 97684
rect 106411 97672 106445 97684
rect 106965 97672 106999 97684
rect 107519 97672 107553 97684
rect 108073 97672 108107 97684
rect 108627 97672 108661 97684
rect 109181 97672 109215 97684
rect 109735 97672 109769 97684
rect 110289 97672 110323 97684
rect 120888 97638 120938 98238
rect 121038 97638 121094 98238
rect 121194 97638 121244 98238
rect 121456 97607 121506 98207
rect 121606 97607 121734 98207
rect 121762 97607 121890 98207
rect 121918 97607 122046 98207
rect 122074 97607 122124 98207
rect 122190 97607 122240 98207
rect 122340 97607 122468 98207
rect 122496 97607 122624 98207
rect 122652 97607 122780 98207
rect 122808 97607 122864 98207
rect 122964 97607 123092 98207
rect 123120 97607 123248 98207
rect 123276 97607 123404 98207
rect 123432 97607 123488 98207
rect 123588 97607 123644 98207
rect 123744 97607 123800 98207
rect 123900 97607 123950 98207
rect 124016 97607 124066 98207
rect 124166 97607 124294 98207
rect 124322 97607 124378 98207
rect 124478 97607 124606 98207
rect 124634 97607 124684 98207
rect 127617 98115 128617 98165
rect 128680 98115 128730 98226
rect 128677 97995 128730 98115
rect 127617 97945 128617 97995
rect 40797 96532 40798 96556
rect 40878 96532 40879 96556
rect 41351 96532 41352 96556
rect 41432 96532 41433 96556
rect 41905 96532 41906 96556
rect 41986 96532 41987 96556
rect 42459 96532 42460 96556
rect 42540 96532 42541 96556
rect 43013 96532 43014 96556
rect 43094 96532 43095 96556
rect 43567 96532 43568 96556
rect 43648 96532 43649 96556
rect 44121 96532 44122 96556
rect 44202 96532 44203 96556
rect 44675 96532 44676 96556
rect 44756 96532 44757 96556
rect 45229 96532 45230 96556
rect 45310 96532 45311 96556
rect 45783 96532 45784 96556
rect 45864 96532 45865 96556
rect 46337 96532 46338 96556
rect 46418 96532 46419 96556
rect 46891 96532 46892 96556
rect 46972 96532 46973 96556
rect 47445 96532 47446 96556
rect 47526 96532 47527 96556
rect 47999 96532 48000 96556
rect 48080 96532 48081 96556
rect 48553 96532 48554 96556
rect 48634 96532 48635 96556
rect 49107 96532 49108 96556
rect 49188 96532 49189 96556
rect 49661 96532 49662 96556
rect 49742 96532 49743 96556
rect 50215 96532 50216 96556
rect 50296 96532 50297 96556
rect 50769 96532 50770 96556
rect 50850 96532 50851 96556
rect 51323 96532 51324 96556
rect 51404 96532 51405 96556
rect 40821 96508 40855 96520
rect 41375 96508 41409 96520
rect 41929 96508 41963 96520
rect 42483 96508 42517 96520
rect 43037 96508 43071 96520
rect 43591 96508 43625 96520
rect 44145 96508 44179 96520
rect 44699 96508 44733 96520
rect 45253 96508 45287 96520
rect 45807 96508 45841 96520
rect 46361 96508 46395 96520
rect 46915 96508 46949 96520
rect 47469 96508 47503 96520
rect 48023 96508 48057 96520
rect 48577 96508 48611 96520
rect 49131 96508 49165 96520
rect 49685 96508 49719 96520
rect 50239 96508 50273 96520
rect 50793 96508 50827 96520
rect 51347 96508 51381 96520
rect -820 95764 -754 95780
rect 6411 95594 6497 95630
rect 3043 95400 3395 95426
rect 3867 95400 4219 95426
rect 4691 95400 5043 95426
rect 5515 95400 5867 95426
rect 3069 92401 3070 95400
rect 3369 92401 3395 95400
rect 3069 92400 3395 92401
rect 3893 92401 3894 95400
rect 4193 92401 4219 95400
rect 3893 92400 4219 92401
rect 4717 92401 4718 95400
rect 5017 92401 5043 95400
rect 4717 92400 5043 92401
rect 5541 92401 5542 95400
rect 5841 92401 5867 95400
rect 5541 92400 5867 92401
rect 6411 92206 6447 95594
rect 6461 92206 6497 95594
rect 7041 95400 7393 95426
rect 7865 95400 8217 95426
rect 8689 95400 9041 95426
rect 9513 95400 9865 95426
rect 7067 92401 7068 95400
rect 7367 92401 7393 95400
rect 7067 92400 7393 92401
rect 7891 92401 7892 95400
rect 8191 92401 8217 95400
rect 7891 92400 8217 92401
rect 8715 92401 8716 95400
rect 9015 92401 9041 95400
rect 8715 92400 9041 92401
rect 9539 92401 9540 95400
rect 9839 92401 9865 95400
rect 22591 95249 22641 96249
rect 23441 95249 23491 96249
rect 23743 95249 23793 96249
rect 25393 95249 25443 96249
rect 25695 95249 25745 96249
rect 27345 95249 27395 96249
rect 27647 95249 27697 96249
rect 29297 95249 29347 96249
rect 29599 95249 29649 96249
rect 31249 95249 31299 96249
rect 31551 95249 31601 96249
rect 33201 95249 33251 96249
rect 68039 95357 68089 96357
rect 68889 95357 68939 96357
rect 69191 95357 69241 96357
rect 70041 95357 70091 96357
rect 88591 96327 88641 97327
rect 89441 96327 89491 97327
rect 89743 96327 89793 97327
rect 90593 96327 90643 97327
rect 127580 97225 127630 97825
rect 127750 97225 127806 97825
rect 127926 97225 127976 97825
rect 128196 97226 128246 97826
rect 128366 97226 128422 97826
rect 128542 97226 128592 97826
rect 128680 97226 128730 97995
rect 128850 97226 128900 98226
rect 128963 98115 129563 98165
rect 128963 98015 128975 98115
rect 130862 98045 130912 98645
rect 131032 98045 131088 98645
rect 131208 98045 131336 98645
rect 131384 98045 131440 98645
rect 131560 98045 131616 98645
rect 131736 98045 131792 98645
rect 131912 98045 132040 98645
rect 132088 98045 132138 98645
rect 128963 97965 129563 98015
rect 128979 97226 129029 97826
rect 129149 97226 129205 97826
rect 129325 97226 129375 97826
rect 129666 97226 129716 97826
rect 129836 97226 129964 97826
rect 130012 97226 130068 97826
rect 130188 97226 130316 97826
rect 130364 97226 130414 97826
rect 130786 97290 130836 97890
rect 130956 97290 131084 97890
rect 131132 97290 131260 97890
rect 131308 97290 131436 97890
rect 131484 97290 131612 97890
rect 131660 97290 131716 97890
rect 131836 97290 131964 97890
rect 132012 97290 132062 97890
rect 123463 97102 123513 97183
rect 119796 96771 119811 96786
rect 119760 96741 119811 96771
rect 119796 96726 119811 96741
rect 120654 96430 120704 97030
rect 120824 96430 120952 97030
rect 121000 96430 121056 97030
rect 121176 96601 121226 97030
rect 121289 96830 121301 97030
rect 123460 96830 123513 97102
rect 121176 96529 121229 96601
rect 123463 96583 123513 96830
rect 123613 96583 123663 97183
rect 123729 96583 123779 97183
rect 123879 96583 124007 97183
rect 124035 96583 124163 97183
rect 124191 96583 124319 97183
rect 124397 96583 124450 97183
rect 121176 96430 121226 96529
rect 121289 96430 121301 96529
rect 123800 96245 124290 96246
rect 124400 96183 124450 96583
rect 124550 96183 124678 97183
rect 124706 96183 124756 97183
rect 124957 96998 124967 97032
rect 124957 96930 124967 96964
rect 124957 96862 124967 96896
rect 124957 96794 124967 96828
rect 124957 96719 124967 96753
rect 124957 96651 124967 96685
rect 124957 96583 124967 96617
rect 124957 96515 124967 96549
rect 124957 96447 124967 96481
rect 124957 96379 124967 96413
rect 124957 96311 124967 96345
rect 124957 96243 124967 96277
rect 124957 96175 124967 96209
rect 97096 96152 97162 96168
rect 124957 96107 124967 96141
rect 22591 94005 22641 95005
rect 23441 94005 23491 95005
rect 23743 94005 23793 95005
rect 25393 94005 25443 95005
rect 25695 94005 25745 95005
rect 27345 94005 27395 95005
rect 27647 94005 27697 95005
rect 29297 94005 29347 95005
rect 29599 94005 29649 95005
rect 31249 94005 31299 95005
rect 31551 94005 31601 95005
rect 33201 94005 33251 95005
rect 38154 94988 38220 95004
rect 45385 94818 45471 94854
rect 42017 94624 42369 94650
rect 42841 94624 43193 94650
rect 43665 94624 44017 94650
rect 44489 94624 44841 94650
rect 22591 92761 22641 93761
rect 23441 92761 23491 93761
rect 23743 92761 23793 93761
rect 25393 92761 25443 93761
rect 25695 92761 25745 93761
rect 27345 92761 27395 93761
rect 27647 92761 27697 93761
rect 29297 92761 29347 93761
rect 29599 92761 29649 93761
rect 31249 92761 31299 93761
rect 31551 92761 31601 93761
rect 33201 92761 33251 93761
rect 9539 92400 9865 92401
rect 6411 92170 6497 92206
rect 42043 91625 42044 94624
rect 42343 91625 42369 94624
rect 42043 91624 42369 91625
rect 42867 91625 42868 94624
rect 43167 91625 43193 94624
rect 42867 91624 43193 91625
rect 43691 91625 43692 94624
rect 43991 91625 44017 94624
rect 43691 91624 44017 91625
rect 44515 91625 44516 94624
rect 44815 91625 44841 94624
rect 44515 91624 44841 91625
rect 45385 91430 45421 94818
rect 45435 91430 45471 94818
rect 46015 94624 46367 94650
rect 46839 94624 47191 94650
rect 47663 94624 48015 94650
rect 48487 94624 48839 94650
rect 46041 91625 46042 94624
rect 46341 91625 46367 94624
rect 46041 91624 46367 91625
rect 46865 91625 46866 94624
rect 47165 91625 47191 94624
rect 46865 91624 47191 91625
rect 47689 91625 47690 94624
rect 47989 91625 48015 94624
rect 47689 91624 48015 91625
rect 48513 91625 48514 94624
rect 48813 91625 48839 94624
rect 59431 94113 59481 95113
rect 60281 94113 60331 95113
rect 60583 94113 60633 95113
rect 62233 94113 62283 95113
rect 62535 94113 62585 95113
rect 64185 94113 64235 95113
rect 64487 94113 64537 95113
rect 66137 94113 66187 95113
rect 66439 94113 66489 95113
rect 68089 94113 68139 95113
rect 68391 94113 68441 95113
rect 70041 94113 70091 95113
rect 79983 95083 80033 96083
rect 80833 95083 80883 96083
rect 81135 95083 81185 96083
rect 82785 95083 82835 96083
rect 83087 95083 83137 96083
rect 84737 95083 84787 96083
rect 85039 95083 85089 96083
rect 86689 95083 86739 96083
rect 86991 95083 87041 96083
rect 88641 95083 88691 96083
rect 88943 95083 88993 96083
rect 90593 95083 90643 96083
rect 125026 96062 125076 97062
rect 125196 96062 125324 97062
rect 125372 96062 125500 97062
rect 125548 96062 125604 97062
rect 125724 96062 125774 97062
rect 125873 96942 125939 96958
rect 126359 96942 126425 96958
rect 125873 96158 125939 96174
rect 126035 96158 126101 96174
rect 126197 96158 126263 96174
rect 126359 96158 126425 96174
rect 126524 96062 126574 97062
rect 126694 96062 126750 97062
rect 126870 96062 126998 97062
rect 127046 96062 127174 97062
rect 127222 96062 127272 97062
rect 127365 96998 127375 97032
rect 127365 96930 127375 96964
rect 127365 96862 127375 96896
rect 127365 96794 127375 96828
rect 127365 96719 127375 96753
rect 127365 96651 127375 96685
rect 127365 96583 127375 96617
rect 127365 96515 127375 96549
rect 127365 96447 127375 96481
rect 127365 96379 127375 96413
rect 127365 96311 127375 96345
rect 127365 96243 127375 96277
rect 127365 96175 127375 96209
rect 127365 96107 127375 96141
rect 127424 96062 127474 97062
rect 127594 96062 127722 97062
rect 127770 96062 127826 97062
rect 127946 96062 127996 97062
rect 128162 96462 128212 97062
rect 128332 96462 128388 97062
rect 128508 96462 128636 97062
rect 128684 96462 128734 97062
rect 128886 96462 128936 97062
rect 129036 96462 129164 97062
rect 129192 96462 129248 97062
rect 129348 96462 129476 97062
rect 129504 96462 129554 97062
rect 129758 96462 129808 97062
rect 129908 96462 130036 97062
rect 130064 96462 130192 97062
rect 130220 96462 130276 97062
rect 130376 96462 130426 97062
rect 132211 96933 132261 96988
rect 104327 95982 104413 96018
rect 100959 95788 101311 95814
rect 101783 95788 102135 95814
rect 102607 95788 102959 95814
rect 103431 95788 103783 95814
rect 59431 92869 59481 93869
rect 60281 92869 60331 93869
rect 60583 92869 60633 93869
rect 62233 92869 62283 93869
rect 62535 92869 62585 93869
rect 64185 92869 64235 93869
rect 64487 92869 64537 93869
rect 66137 92869 66187 93869
rect 66439 92869 66489 93869
rect 68089 92869 68139 93869
rect 68391 92869 68441 93869
rect 70041 92869 70091 93869
rect 79983 93839 80033 94839
rect 80833 93839 80883 94839
rect 81135 93839 81185 94839
rect 82785 93839 82835 94839
rect 83087 93839 83137 94839
rect 84737 93839 84787 94839
rect 85039 93839 85089 94839
rect 86689 93839 86739 94839
rect 86991 93839 87041 94839
rect 88641 93839 88691 94839
rect 88943 93839 88993 94839
rect 90593 93839 90643 94839
rect 59431 91625 59481 92625
rect 60281 91625 60331 92625
rect 60583 91625 60633 92625
rect 62233 91625 62283 92625
rect 62535 91625 62585 92625
rect 64185 91625 64235 92625
rect 64487 91625 64537 92625
rect 66137 91625 66187 92625
rect 66439 91625 66489 92625
rect 68089 91625 68139 92625
rect 68391 91625 68441 92625
rect 70041 91625 70091 92625
rect 79983 92595 80033 93595
rect 80833 92595 80883 93595
rect 81135 92595 81185 93595
rect 82785 92595 82835 93595
rect 83087 92595 83137 93595
rect 84737 92595 84787 93595
rect 85039 92595 85089 93595
rect 86689 92595 86739 93595
rect 86991 92595 87041 93595
rect 88641 92595 88691 93595
rect 88943 92595 88993 93595
rect 90593 92595 90643 93595
rect 100985 92789 100986 95788
rect 101285 92789 101311 95788
rect 100985 92788 101311 92789
rect 101809 92789 101810 95788
rect 102109 92789 102135 95788
rect 101809 92788 102135 92789
rect 102633 92789 102634 95788
rect 102933 92789 102959 95788
rect 102633 92788 102959 92789
rect 103457 92789 103458 95788
rect 103757 92789 103783 95788
rect 103457 92788 103783 92789
rect 104327 92594 104363 95982
rect 104377 92594 104413 95982
rect 104957 95788 105309 95814
rect 105781 95788 106133 95814
rect 106605 95788 106957 95814
rect 107429 95788 107781 95814
rect 104983 92789 104984 95788
rect 105283 92789 105309 95788
rect 104983 92788 105309 92789
rect 105807 92789 105808 95788
rect 106107 92789 106133 95788
rect 105807 92788 106133 92789
rect 106631 92789 106632 95788
rect 106931 92789 106957 95788
rect 106631 92788 106957 92789
rect 107455 92789 107456 95788
rect 107755 92789 107781 95788
rect 119826 95382 119879 95532
rect 119829 94932 119879 95382
rect 119999 94932 120055 95532
rect 120175 94932 120231 95532
rect 120351 94932 120407 95532
rect 120527 94932 120577 95532
rect 120643 94932 120693 95532
rect 120813 94932 120869 95532
rect 120989 94932 121045 95532
rect 121165 94932 121215 95532
rect 121486 95332 121666 95532
rect 121722 95332 121902 95532
rect 123456 95332 123636 95532
rect 123692 95332 123872 95532
rect 121722 95197 121902 95234
rect 123456 95197 123636 95234
rect 124143 94932 124193 95532
rect 124313 94932 124369 95532
rect 124489 94932 124545 95532
rect 124665 94932 124715 95532
rect 124797 94932 124847 95532
rect 124967 94932 125023 95532
rect 125143 94932 125199 95532
rect 125319 94932 125369 95532
rect 125640 95332 125820 95532
rect 125876 95332 126056 95532
rect 127610 95332 127790 95532
rect 127846 95332 128026 95532
rect 125876 95197 126056 95234
rect 127610 95197 127790 95234
rect 128297 94932 128347 95532
rect 128467 94932 128523 95532
rect 128643 94932 128699 95532
rect 128819 94932 128869 95532
rect 128951 94932 129001 95532
rect 129121 94932 129177 95532
rect 129297 94932 129353 95532
rect 129473 94932 129523 95532
rect 129794 95332 129974 95532
rect 130030 95332 130210 95532
rect 131764 95332 131944 95532
rect 132000 95332 132180 95532
rect 130030 95197 130210 95234
rect 131764 95197 131944 95234
rect 132451 94932 132501 95532
rect 132621 94932 132677 95532
rect 132797 94932 132853 95532
rect 132973 94932 133023 95532
rect 133204 94534 133228 94558
rect 133625 94534 133649 94558
rect 133228 94510 133252 94525
rect 133601 94510 133625 94525
rect 133032 94354 133056 94378
rect 133057 94330 133080 94354
rect 119452 93516 119502 94116
rect 119622 93516 119678 94116
rect 119798 93516 119848 94116
rect 121341 93724 121391 94324
rect 121511 93724 121561 94324
rect 121937 93719 121987 94319
rect 122107 93719 122163 94319
rect 122283 94072 122333 94319
rect 122396 94169 122408 94319
rect 123022 94169 123075 94319
rect 123025 94072 123075 94169
rect 122283 94000 122336 94072
rect 122283 93719 122333 94000
rect 122396 93850 122408 94000
rect 123022 93850 123075 94072
rect 123025 93719 123075 93850
rect 123195 93719 123251 94319
rect 123371 93719 123421 94319
rect 123797 93724 123847 94324
rect 123967 93724 124017 94324
rect 125495 93724 125545 94324
rect 125665 93724 125715 94324
rect 126091 93719 126141 94319
rect 126261 93719 126317 94319
rect 126437 94072 126487 94319
rect 126550 94169 126562 94319
rect 127176 94169 127229 94319
rect 127179 94072 127229 94169
rect 126437 94000 126490 94072
rect 126437 93719 126487 94000
rect 126550 93850 126562 94000
rect 127176 93850 127229 94072
rect 127179 93719 127229 93850
rect 127349 93719 127405 94319
rect 127525 93719 127575 94319
rect 127951 93724 128001 94324
rect 128121 93724 128171 94324
rect 129649 93724 129699 94324
rect 129819 93724 129869 94324
rect 130245 93719 130295 94319
rect 130415 93719 130471 94319
rect 130591 94072 130641 94319
rect 130704 94169 130716 94319
rect 131330 94169 131383 94319
rect 131333 94072 131383 94169
rect 130591 94000 130644 94072
rect 130591 93719 130641 94000
rect 130704 93850 130716 94000
rect 131330 93850 131383 94072
rect 131333 93719 131383 93850
rect 131503 93719 131559 94319
rect 131679 93719 131729 94319
rect 132105 93724 132155 94324
rect 132275 93724 132325 94324
rect 133252 94266 133286 94290
rect 133322 94266 133356 94290
rect 133392 94266 133426 94290
rect 133462 94266 133496 94290
rect 133532 94266 133566 94290
rect 133602 94266 133625 94290
rect 133057 94232 133080 94256
rect 133032 94208 133056 94232
rect 120880 93397 120914 93421
rect 120948 93397 120982 93421
rect 121016 93397 121050 93421
rect 121084 93397 121118 93421
rect 121152 93397 121186 93421
rect 121220 93397 121254 93421
rect 121288 93397 121322 93421
rect 121356 93397 121390 93421
rect 121424 93397 121458 93421
rect 121492 93397 121526 93421
rect 121560 93397 121594 93421
rect 121628 93397 121662 93421
rect 121696 93397 121730 93421
rect 121764 93397 121798 93421
rect 121832 93397 121866 93421
rect 121900 93397 121934 93421
rect 121968 93397 122002 93421
rect 122036 93397 122070 93421
rect 122104 93397 122138 93421
rect 122172 93397 122206 93421
rect 122240 93397 122274 93421
rect 122308 93397 122342 93421
rect 122376 93397 122410 93421
rect 122444 93397 122478 93421
rect 122512 93397 122546 93421
rect 122580 93397 122614 93421
rect 122648 93397 122682 93421
rect 122716 93397 122750 93421
rect 122784 93397 122818 93421
rect 122852 93397 122886 93421
rect 122920 93397 122954 93421
rect 122988 93397 123022 93421
rect 123056 93397 123090 93421
rect 123124 93397 123158 93421
rect 123192 93397 123226 93421
rect 123260 93397 123294 93421
rect 123328 93397 123362 93421
rect 123396 93397 123430 93421
rect 123464 93397 123498 93421
rect 123532 93397 123566 93421
rect 123600 93397 123634 93421
rect 123668 93397 123702 93421
rect 123736 93397 123770 93421
rect 123804 93397 123838 93421
rect 123872 93397 123906 93421
rect 123940 93397 123974 93421
rect 124008 93397 124042 93421
rect 124076 93397 124110 93421
rect 124144 93397 124178 93421
rect 124212 93397 124246 93421
rect 124280 93397 124314 93421
rect 124348 93397 124382 93421
rect 124416 93397 124450 93421
rect 124484 93397 124518 93421
rect 124552 93397 124586 93421
rect 124620 93397 124654 93421
rect 124688 93397 124722 93421
rect 124756 93397 124790 93421
rect 124824 93397 124858 93421
rect 124892 93397 124926 93421
rect 124960 93397 124994 93421
rect 125028 93397 125062 93421
rect 125096 93397 125130 93421
rect 125164 93397 125198 93421
rect 125232 93397 125266 93421
rect 125300 93397 125334 93421
rect 125368 93397 125402 93421
rect 125436 93397 125470 93421
rect 125504 93397 125538 93421
rect 125572 93397 125606 93421
rect 125640 93397 125674 93421
rect 125708 93397 125742 93421
rect 125776 93397 125810 93421
rect 125844 93397 125878 93421
rect 125912 93397 125946 93421
rect 125980 93397 126014 93421
rect 126048 93397 126082 93421
rect 126116 93397 126150 93421
rect 126184 93397 126218 93421
rect 126252 93397 126286 93421
rect 126320 93397 126354 93421
rect 126388 93397 126422 93421
rect 126456 93397 126490 93421
rect 126524 93397 126558 93421
rect 126592 93397 126626 93421
rect 126660 93397 126694 93421
rect 126728 93397 126762 93421
rect 126796 93397 126830 93421
rect 126864 93397 126898 93421
rect 126932 93397 126966 93421
rect 127000 93397 127034 93421
rect 127068 93397 127102 93421
rect 127136 93397 127170 93421
rect 127204 93397 127238 93421
rect 127272 93397 127306 93421
rect 127340 93397 127374 93421
rect 127408 93397 127442 93421
rect 127476 93397 127510 93421
rect 127544 93397 127578 93421
rect 127612 93397 127646 93421
rect 127680 93397 127714 93421
rect 127748 93397 127782 93421
rect 127816 93397 127850 93421
rect 127884 93397 127918 93421
rect 127952 93397 127986 93421
rect 128020 93397 128054 93421
rect 128088 93397 128122 93421
rect 128156 93397 128190 93421
rect 128224 93397 128258 93421
rect 128358 93397 128392 93421
rect 128426 93397 128460 93421
rect 128494 93397 128528 93421
rect 128562 93397 128596 93421
rect 128630 93397 128664 93421
rect 128698 93397 128732 93421
rect 128766 93397 128800 93421
rect 128834 93397 128868 93421
rect 128902 93397 128936 93421
rect 128970 93397 129004 93421
rect 129038 93397 129072 93421
rect 129106 93397 129140 93421
rect 129174 93397 129208 93421
rect 129242 93397 129276 93421
rect 129310 93397 129344 93421
rect 129378 93397 129412 93421
rect 129446 93397 129480 93421
rect 129514 93397 129548 93421
rect 129582 93397 129616 93421
rect 129650 93397 129684 93421
rect 129718 93397 129752 93421
rect 129786 93397 129820 93421
rect 129854 93397 129888 93421
rect 129922 93397 129956 93421
rect 129990 93397 130024 93421
rect 130058 93397 130092 93421
rect 130126 93397 130160 93421
rect 130194 93397 130228 93421
rect 130262 93397 130296 93421
rect 130330 93397 130364 93421
rect 130398 93397 130432 93421
rect 130466 93397 130500 93421
rect 130534 93397 130568 93421
rect 130602 93397 130636 93421
rect 130670 93397 130704 93421
rect 130738 93397 130772 93421
rect 130806 93397 130840 93421
rect 130874 93397 130908 93421
rect 130942 93397 130976 93421
rect 131010 93397 131044 93421
rect 131078 93397 131112 93421
rect 131146 93397 131180 93421
rect 131214 93397 131248 93421
rect 131282 93397 131316 93421
rect 131350 93397 131384 93421
rect 131418 93397 131452 93421
rect 128334 93363 128362 93397
rect 107455 92788 107781 92789
rect 104327 92558 104413 92594
rect 48513 91624 48839 91625
rect 45385 91394 45471 91430
rect 1188 85320 1254 85336
rect 2211 83550 2212 83574
rect 2292 83550 2293 83574
rect 2765 83550 2766 83574
rect 2846 83550 2847 83574
rect 3319 83550 3320 83574
rect 3400 83550 3401 83574
rect 3873 83550 3874 83574
rect 3954 83550 3955 83574
rect 4427 83550 4428 83574
rect 4508 83550 4509 83574
rect 4981 83550 4982 83574
rect 5062 83550 5063 83574
rect 5535 83550 5536 83574
rect 5616 83550 5617 83574
rect 6089 83550 6090 83574
rect 6170 83550 6171 83574
rect 6643 83550 6644 83574
rect 6724 83550 6725 83574
rect 7197 83550 7198 83574
rect 7278 83550 7279 83574
rect 7751 83550 7752 83574
rect 7832 83550 7833 83574
rect 8305 83550 8306 83574
rect 8386 83550 8387 83574
rect 8859 83550 8860 83574
rect 8940 83550 8941 83574
rect 9413 83550 9414 83574
rect 9494 83550 9495 83574
rect 9967 83550 9968 83574
rect 10048 83550 10049 83574
rect 10521 83550 10522 83574
rect 10602 83550 10603 83574
rect 11075 83550 11076 83574
rect 11156 83550 11157 83574
rect 11629 83550 11630 83574
rect 11710 83550 11711 83574
rect 12183 83550 12184 83574
rect 12264 83550 12265 83574
rect 12737 83550 12738 83574
rect 12818 83550 12819 83574
rect 2235 83526 2269 83538
rect 2789 83526 2823 83538
rect 3343 83526 3377 83538
rect 3897 83526 3931 83538
rect 4451 83526 4485 83538
rect 5005 83526 5039 83538
rect 5559 83526 5593 83538
rect 6113 83526 6147 83538
rect 6667 83526 6701 83538
rect 7221 83526 7255 83538
rect 7775 83526 7809 83538
rect 8329 83526 8363 83538
rect 8883 83526 8917 83538
rect 9437 83526 9471 83538
rect 9991 83526 10025 83538
rect 10545 83526 10579 83538
rect 11099 83526 11133 83538
rect 11653 83526 11687 83538
rect 12207 83526 12241 83538
rect 12761 83526 12795 83538
rect 21232 83370 21304 85370
rect 21503 83403 21621 85297
rect 21892 83370 21952 85370
rect 22152 83370 22224 85370
rect 22423 83403 22541 85297
rect 22812 83370 22872 85370
rect 23072 83370 23144 85370
rect 23343 83403 23461 85297
rect 23732 83370 23792 85370
rect 23992 83370 24064 85370
rect 24263 83403 24381 85297
rect 24652 83370 24712 85370
rect 24912 83370 24984 85370
rect 25183 83403 25301 85297
rect 25572 83370 25632 85370
rect 25832 83370 25904 85370
rect 26103 83403 26221 85297
rect 26492 83370 26552 85370
rect 26752 83370 26824 85370
rect 27023 83403 27141 85297
rect 27412 83370 27472 85370
rect 27672 83370 27744 85370
rect 27943 83403 28061 85297
rect 28332 83370 28392 85370
rect 28592 83370 28664 85370
rect 28863 83403 28981 85297
rect 29252 83370 29312 85370
rect 29512 83370 29584 85370
rect 29783 83403 29901 85297
rect 30172 83370 30232 85370
rect 30432 83370 30504 85370
rect 30703 83403 30821 85297
rect 31092 83370 31152 85370
rect 41010 83564 41082 85564
rect 41281 83597 41399 85491
rect 41670 83564 41730 85564
rect 41930 83564 42002 85564
rect 42201 83597 42319 85491
rect 42590 83564 42650 85564
rect 42850 83564 42922 85564
rect 43121 83597 43239 85491
rect 43510 83564 43570 85564
rect 43770 83564 43842 85564
rect 44041 83597 44159 85491
rect 44430 83564 44490 85564
rect 44690 83564 44762 85564
rect 44961 83597 45079 85491
rect 45350 83564 45410 85564
rect 45610 83564 45682 85564
rect 45881 83597 45999 85491
rect 46270 83564 46330 85564
rect 46530 83564 46602 85564
rect 46801 83597 46919 85491
rect 47190 83564 47250 85564
rect 47450 83564 47522 85564
rect 47721 83597 47839 85491
rect 48110 83564 48170 85564
rect 48370 83564 48442 85564
rect 48641 83597 48759 85491
rect 49030 83564 49090 85564
rect 49290 83564 49362 85564
rect 49561 83597 49679 85491
rect 49950 83564 50010 85564
rect 50210 83564 50282 85564
rect 50481 83597 50599 85491
rect 50870 83564 50930 85564
rect 61684 83574 61750 83590
rect 80686 83380 80752 83396
rect 2765 81550 2766 81574
rect 2846 81550 2847 81574
rect 3319 81550 3320 81574
rect 3400 81550 3401 81574
rect 3873 81550 3874 81574
rect 3954 81550 3955 81574
rect 4427 81550 4428 81574
rect 4508 81550 4509 81574
rect 4981 81550 4982 81574
rect 5062 81550 5063 81574
rect 5535 81550 5536 81574
rect 5616 81550 5617 81574
rect 6089 81550 6090 81574
rect 6170 81550 6171 81574
rect 6643 81550 6644 81574
rect 6724 81550 6725 81574
rect 7197 81550 7198 81574
rect 7278 81550 7279 81574
rect 7751 81550 7752 81574
rect 7832 81550 7833 81574
rect 8305 81550 8306 81574
rect 8386 81550 8387 81574
rect 8859 81550 8860 81574
rect 8940 81550 8941 81574
rect 9413 81550 9414 81574
rect 9494 81550 9495 81574
rect 9967 81550 9968 81574
rect 10048 81550 10049 81574
rect 10521 81550 10522 81574
rect 10602 81550 10603 81574
rect 11075 81550 11076 81574
rect 11156 81550 11157 81574
rect 11629 81550 11630 81574
rect 11710 81550 11711 81574
rect 12183 81550 12184 81574
rect 12264 81550 12265 81574
rect 12737 81550 12738 81574
rect 12818 81550 12819 81574
rect 2789 81526 2823 81538
rect 3343 81526 3377 81538
rect 3897 81526 3931 81538
rect 4451 81526 4485 81538
rect 5005 81526 5039 81538
rect 5559 81526 5593 81538
rect 6113 81526 6147 81538
rect 6667 81526 6701 81538
rect 7221 81526 7255 81538
rect 7775 81526 7809 81538
rect 8329 81526 8363 81538
rect 8883 81526 8917 81538
rect 9437 81526 9471 81538
rect 9991 81526 10025 81538
rect 10545 81526 10579 81538
rect 11099 81526 11133 81538
rect 11653 81526 11687 81538
rect 12207 81526 12241 81538
rect 12761 81526 12795 81538
rect 2705 79550 2706 79574
rect 2786 79550 2787 79574
rect 3541 79550 3542 79574
rect 3622 79550 3623 79574
rect 4377 79550 4378 79574
rect 4458 79550 4459 79574
rect 5213 79550 5214 79574
rect 5294 79550 5295 79574
rect 6049 79550 6050 79574
rect 6130 79550 6131 79574
rect 6885 79550 6886 79574
rect 6966 79550 6967 79574
rect 7721 79550 7722 79574
rect 7802 79550 7803 79574
rect 8557 79550 8558 79574
rect 8638 79550 8639 79574
rect 9393 79550 9394 79574
rect 9474 79550 9475 79574
rect 10229 79550 10230 79574
rect 10310 79550 10311 79574
rect 11065 79550 11066 79574
rect 11146 79550 11147 79574
rect 11901 79550 11902 79574
rect 11982 79550 11983 79574
rect 12737 79550 12738 79574
rect 12818 79550 12819 79574
rect 2729 79526 2763 79538
rect 3565 79526 3599 79538
rect 4401 79526 4435 79538
rect 5237 79526 5271 79538
rect 6073 79526 6107 79538
rect 6909 79526 6943 79538
rect 7745 79526 7779 79538
rect 8581 79526 8615 79538
rect 9417 79526 9451 79538
rect 10253 79526 10287 79538
rect 11089 79526 11123 79538
rect 11925 79526 11959 79538
rect 12761 79526 12795 79538
rect 21232 78770 21304 82770
rect 21503 78803 21621 82737
rect 21892 78770 21952 82770
rect 22152 78770 22224 82770
rect 22423 78803 22541 82737
rect 22812 78770 22872 82770
rect 23072 78770 23144 82770
rect 23343 78803 23461 82737
rect 23732 78770 23792 82770
rect 23992 78770 24064 82770
rect 24263 78803 24381 82737
rect 24652 78770 24712 82770
rect 24912 78770 24984 82770
rect 25183 78803 25301 82737
rect 25572 78770 25632 82770
rect 25832 78770 25904 82770
rect 26103 78803 26221 82737
rect 26492 78770 26552 82770
rect 26752 78770 26824 82770
rect 27023 78803 27141 82737
rect 27412 78770 27472 82770
rect 27672 78770 27744 82770
rect 27943 78803 28061 82737
rect 28332 78770 28392 82770
rect 28592 78770 28664 82770
rect 28863 78803 28981 82737
rect 29252 78770 29312 82770
rect 29512 78770 29584 82770
rect 29783 78803 29901 82737
rect 30172 78770 30232 82770
rect 30432 78770 30504 82770
rect 30703 78803 30821 82737
rect 31092 78770 31152 82770
rect 41010 78964 41082 82964
rect 41281 78997 41399 82931
rect 41670 78964 41730 82964
rect 41930 78964 42002 82964
rect 42201 78997 42319 82931
rect 42590 78964 42650 82964
rect 42850 78964 42922 82964
rect 43121 78997 43239 82931
rect 43510 78964 43570 82964
rect 43770 78964 43842 82964
rect 44041 78997 44159 82931
rect 44430 78964 44490 82964
rect 44690 78964 44762 82964
rect 44961 78997 45079 82931
rect 45350 78964 45410 82964
rect 45610 78964 45682 82964
rect 45881 78997 45999 82931
rect 46270 78964 46330 82964
rect 46530 78964 46602 82964
rect 46801 78997 46919 82931
rect 47190 78964 47250 82964
rect 47450 78964 47522 82964
rect 47721 78997 47839 82931
rect 48110 78964 48170 82964
rect 48370 78964 48442 82964
rect 48641 78997 48759 82931
rect 49030 78964 49090 82964
rect 49290 78964 49362 82964
rect 49561 78997 49679 82931
rect 49950 78964 50010 82964
rect 50210 78964 50282 82964
rect 50481 78997 50599 82931
rect 50870 78964 50930 82964
rect 62707 81804 62708 81828
rect 62788 81804 62789 81828
rect 63261 81804 63262 81828
rect 63342 81804 63343 81828
rect 63815 81804 63816 81828
rect 63896 81804 63897 81828
rect 64369 81804 64370 81828
rect 64450 81804 64451 81828
rect 64923 81804 64924 81828
rect 65004 81804 65005 81828
rect 65477 81804 65478 81828
rect 65558 81804 65559 81828
rect 66031 81804 66032 81828
rect 66112 81804 66113 81828
rect 66585 81804 66586 81828
rect 66666 81804 66667 81828
rect 67139 81804 67140 81828
rect 67220 81804 67221 81828
rect 67693 81804 67694 81828
rect 67774 81804 67775 81828
rect 68247 81804 68248 81828
rect 68328 81804 68329 81828
rect 68801 81804 68802 81828
rect 68882 81804 68883 81828
rect 69355 81804 69356 81828
rect 69436 81804 69437 81828
rect 69909 81804 69910 81828
rect 69990 81804 69991 81828
rect 70463 81804 70464 81828
rect 70544 81804 70545 81828
rect 71017 81804 71018 81828
rect 71098 81804 71099 81828
rect 71571 81804 71572 81828
rect 71652 81804 71653 81828
rect 72125 81804 72126 81828
rect 72206 81804 72207 81828
rect 72679 81804 72680 81828
rect 72760 81804 72761 81828
rect 73233 81804 73234 81828
rect 73314 81804 73315 81828
rect 62731 81780 62765 81792
rect 63285 81780 63319 81792
rect 63839 81780 63873 81792
rect 64393 81780 64427 81792
rect 64947 81780 64981 81792
rect 65501 81780 65535 81792
rect 66055 81780 66089 81792
rect 66609 81780 66643 81792
rect 67163 81780 67197 81792
rect 67717 81780 67751 81792
rect 68271 81780 68305 81792
rect 68825 81780 68859 81792
rect 69379 81780 69413 81792
rect 69933 81780 69967 81792
rect 70487 81780 70521 81792
rect 71041 81780 71075 81792
rect 71595 81780 71629 81792
rect 72149 81780 72183 81792
rect 72703 81780 72737 81792
rect 73257 81780 73291 81792
rect 81709 81610 81710 81634
rect 81790 81610 81791 81634
rect 82263 81610 82264 81634
rect 82344 81610 82345 81634
rect 82817 81610 82818 81634
rect 82898 81610 82899 81634
rect 83371 81610 83372 81634
rect 83452 81610 83453 81634
rect 83925 81610 83926 81634
rect 84006 81610 84007 81634
rect 84479 81610 84480 81634
rect 84560 81610 84561 81634
rect 85033 81610 85034 81634
rect 85114 81610 85115 81634
rect 85587 81610 85588 81634
rect 85668 81610 85669 81634
rect 86141 81610 86142 81634
rect 86222 81610 86223 81634
rect 86695 81610 86696 81634
rect 86776 81610 86777 81634
rect 87249 81610 87250 81634
rect 87330 81610 87331 81634
rect 87803 81610 87804 81634
rect 87884 81610 87885 81634
rect 88357 81610 88358 81634
rect 88438 81610 88439 81634
rect 88911 81610 88912 81634
rect 88992 81610 88993 81634
rect 89465 81610 89466 81634
rect 89546 81610 89547 81634
rect 90019 81610 90020 81634
rect 90100 81610 90101 81634
rect 90573 81610 90574 81634
rect 90654 81610 90655 81634
rect 91127 81610 91128 81634
rect 91208 81610 91209 81634
rect 91681 81610 91682 81634
rect 91762 81610 91763 81634
rect 92235 81610 92236 81634
rect 92316 81610 92317 81634
rect 81733 81586 81767 81598
rect 82287 81586 82321 81598
rect 82841 81586 82875 81598
rect 83395 81586 83429 81598
rect 83949 81586 83983 81598
rect 84503 81586 84537 81598
rect 85057 81586 85091 81598
rect 85611 81586 85645 81598
rect 86165 81586 86199 81598
rect 86719 81586 86753 81598
rect 87273 81586 87307 81598
rect 87827 81586 87861 81598
rect 88381 81586 88415 81598
rect 88935 81586 88969 81598
rect 89489 81586 89523 81598
rect 90043 81586 90077 81598
rect 90597 81586 90631 81598
rect 91151 81586 91185 81598
rect 91705 81586 91739 81598
rect 92259 81586 92293 81598
rect 103638 81596 103710 83596
rect 103909 81629 104027 83523
rect 104298 81596 104358 83596
rect 104558 81596 104630 83596
rect 104829 81629 104947 83523
rect 105218 81596 105278 83596
rect 105478 81596 105550 83596
rect 105749 81629 105867 83523
rect 106138 81596 106198 83596
rect 106398 81596 106470 83596
rect 106669 81629 106787 83523
rect 107058 81596 107118 83596
rect 107318 81596 107390 83596
rect 107589 81629 107707 83523
rect 107978 81596 108038 83596
rect 108238 81596 108310 83596
rect 108509 81629 108627 83523
rect 108898 81596 108958 83596
rect 109158 81596 109230 83596
rect 109429 81629 109547 83523
rect 109818 81596 109878 83596
rect 110078 81596 110150 83596
rect 110349 81629 110467 83523
rect 110738 81596 110798 83596
rect 110998 81596 111070 83596
rect 111269 81629 111387 83523
rect 111658 81596 111718 83596
rect 111918 81596 111990 83596
rect 112189 81629 112307 83523
rect 112578 81596 112638 83596
rect 112838 81596 112910 83596
rect 113109 81629 113227 83523
rect 113498 81596 113558 83596
rect 63261 79804 63262 79828
rect 63342 79804 63343 79828
rect 63815 79804 63816 79828
rect 63896 79804 63897 79828
rect 64369 79804 64370 79828
rect 64450 79804 64451 79828
rect 64923 79804 64924 79828
rect 65004 79804 65005 79828
rect 65477 79804 65478 79828
rect 65558 79804 65559 79828
rect 66031 79804 66032 79828
rect 66112 79804 66113 79828
rect 66585 79804 66586 79828
rect 66666 79804 66667 79828
rect 67139 79804 67140 79828
rect 67220 79804 67221 79828
rect 67693 79804 67694 79828
rect 67774 79804 67775 79828
rect 68247 79804 68248 79828
rect 68328 79804 68329 79828
rect 68801 79804 68802 79828
rect 68882 79804 68883 79828
rect 69355 79804 69356 79828
rect 69436 79804 69437 79828
rect 69909 79804 69910 79828
rect 69990 79804 69991 79828
rect 70463 79804 70464 79828
rect 70544 79804 70545 79828
rect 71017 79804 71018 79828
rect 71098 79804 71099 79828
rect 71571 79804 71572 79828
rect 71652 79804 71653 79828
rect 72125 79804 72126 79828
rect 72206 79804 72207 79828
rect 72679 79804 72680 79828
rect 72760 79804 72761 79828
rect 73233 79804 73234 79828
rect 73314 79804 73315 79828
rect 63285 79780 63319 79792
rect 63839 79780 63873 79792
rect 64393 79780 64427 79792
rect 64947 79780 64981 79792
rect 65501 79780 65535 79792
rect 66055 79780 66089 79792
rect 66609 79780 66643 79792
rect 67163 79780 67197 79792
rect 67717 79780 67751 79792
rect 68271 79780 68305 79792
rect 68825 79780 68859 79792
rect 69379 79780 69413 79792
rect 69933 79780 69967 79792
rect 70487 79780 70521 79792
rect 71041 79780 71075 79792
rect 71595 79780 71629 79792
rect 72149 79780 72183 79792
rect 72703 79780 72737 79792
rect 73257 79780 73291 79792
rect 82263 79610 82264 79634
rect 82344 79610 82345 79634
rect 82817 79610 82818 79634
rect 82898 79610 82899 79634
rect 83371 79610 83372 79634
rect 83452 79610 83453 79634
rect 83925 79610 83926 79634
rect 84006 79610 84007 79634
rect 84479 79610 84480 79634
rect 84560 79610 84561 79634
rect 85033 79610 85034 79634
rect 85114 79610 85115 79634
rect 85587 79610 85588 79634
rect 85668 79610 85669 79634
rect 86141 79610 86142 79634
rect 86222 79610 86223 79634
rect 86695 79610 86696 79634
rect 86776 79610 86777 79634
rect 87249 79610 87250 79634
rect 87330 79610 87331 79634
rect 87803 79610 87804 79634
rect 87884 79610 87885 79634
rect 88357 79610 88358 79634
rect 88438 79610 88439 79634
rect 88911 79610 88912 79634
rect 88992 79610 88993 79634
rect 89465 79610 89466 79634
rect 89546 79610 89547 79634
rect 90019 79610 90020 79634
rect 90100 79610 90101 79634
rect 90573 79610 90574 79634
rect 90654 79610 90655 79634
rect 91127 79610 91128 79634
rect 91208 79610 91209 79634
rect 91681 79610 91682 79634
rect 91762 79610 91763 79634
rect 92235 79610 92236 79634
rect 92316 79610 92317 79634
rect 82287 79586 82321 79598
rect 82841 79586 82875 79598
rect 83395 79586 83429 79598
rect 83949 79586 83983 79598
rect 84503 79586 84537 79598
rect 85057 79586 85091 79598
rect 85611 79586 85645 79598
rect 86165 79586 86199 79598
rect 86719 79586 86753 79598
rect 87273 79586 87307 79598
rect 87827 79586 87861 79598
rect 88381 79586 88415 79598
rect 88935 79586 88969 79598
rect 89489 79586 89523 79598
rect 90043 79586 90077 79598
rect 90597 79586 90631 79598
rect 91151 79586 91185 79598
rect 91705 79586 91739 79598
rect 92259 79586 92293 79598
rect 2705 77550 2706 77574
rect 2786 77550 2787 77574
rect 3541 77550 3542 77574
rect 3622 77550 3623 77574
rect 4377 77550 4378 77574
rect 4458 77550 4459 77574
rect 5213 77550 5214 77574
rect 5294 77550 5295 77574
rect 6049 77550 6050 77574
rect 6130 77550 6131 77574
rect 6885 77550 6886 77574
rect 6966 77550 6967 77574
rect 7721 77550 7722 77574
rect 7802 77550 7803 77574
rect 8557 77550 8558 77574
rect 8638 77550 8639 77574
rect 9393 77550 9394 77574
rect 9474 77550 9475 77574
rect 10229 77550 10230 77574
rect 10310 77550 10311 77574
rect 11065 77550 11066 77574
rect 11146 77550 11147 77574
rect 11901 77550 11902 77574
rect 11982 77550 11983 77574
rect 12737 77550 12738 77574
rect 12818 77550 12819 77574
rect 2729 77526 2763 77538
rect 3565 77526 3599 77538
rect 4401 77526 4435 77538
rect 5237 77526 5271 77538
rect 6073 77526 6107 77538
rect 6909 77526 6943 77538
rect 7745 77526 7779 77538
rect 8581 77526 8615 77538
rect 9417 77526 9451 77538
rect 10253 77526 10287 77538
rect 11089 77526 11123 77538
rect 11925 77526 11959 77538
rect 12761 77526 12795 77538
rect 2705 75550 2706 75574
rect 2786 75550 2787 75574
rect 3541 75550 3542 75574
rect 3622 75550 3623 75574
rect 4377 75550 4378 75574
rect 4458 75550 4459 75574
rect 5213 75550 5214 75574
rect 5294 75550 5295 75574
rect 6049 75550 6050 75574
rect 6130 75550 6131 75574
rect 6885 75550 6886 75574
rect 6966 75550 6967 75574
rect 7721 75550 7722 75574
rect 7802 75550 7803 75574
rect 8557 75550 8558 75574
rect 8638 75550 8639 75574
rect 9393 75550 9394 75574
rect 9474 75550 9475 75574
rect 10229 75550 10230 75574
rect 10310 75550 10311 75574
rect 11065 75550 11066 75574
rect 11146 75550 11147 75574
rect 11901 75550 11902 75574
rect 11982 75550 11983 75574
rect 12737 75550 12738 75574
rect 12818 75550 12819 75574
rect 2729 75526 2763 75538
rect 3565 75526 3599 75538
rect 4401 75526 4435 75538
rect 5237 75526 5271 75538
rect 6073 75526 6107 75538
rect 6909 75526 6943 75538
rect 7745 75526 7779 75538
rect 8581 75526 8615 75538
rect 9417 75526 9451 75538
rect 10253 75526 10287 75538
rect 11089 75526 11123 75538
rect 11925 75526 11959 75538
rect 12761 75526 12795 75538
rect 21232 74170 21304 78170
rect 21503 74203 21621 78137
rect 21892 74170 21952 78170
rect 22152 74170 22224 78170
rect 22423 74203 22541 78137
rect 22812 74170 22872 78170
rect 23072 74170 23144 78170
rect 23343 74203 23461 78137
rect 23732 74170 23792 78170
rect 23992 74170 24064 78170
rect 24263 74203 24381 78137
rect 24652 74170 24712 78170
rect 24912 74170 24984 78170
rect 25183 74203 25301 78137
rect 25572 74170 25632 78170
rect 25832 74170 25904 78170
rect 26103 74203 26221 78137
rect 26492 74170 26552 78170
rect 26752 74170 26824 78170
rect 27023 74203 27141 78137
rect 27412 74170 27472 78170
rect 27672 74170 27744 78170
rect 27943 74203 28061 78137
rect 28332 74170 28392 78170
rect 28592 74170 28664 78170
rect 28863 74203 28981 78137
rect 29252 74170 29312 78170
rect 29512 74170 29584 78170
rect 29783 74203 29901 78137
rect 30172 74170 30232 78170
rect 30432 74170 30504 78170
rect 30703 74203 30821 78137
rect 31092 74170 31152 78170
rect 41010 74364 41082 78364
rect 41281 74397 41399 78331
rect 41670 74364 41730 78364
rect 41930 74364 42002 78364
rect 42201 74397 42319 78331
rect 42590 74364 42650 78364
rect 42850 74364 42922 78364
rect 43121 74397 43239 78331
rect 43510 74364 43570 78364
rect 43770 74364 43842 78364
rect 44041 74397 44159 78331
rect 44430 74364 44490 78364
rect 44690 74364 44762 78364
rect 44961 74397 45079 78331
rect 45350 74364 45410 78364
rect 45610 74364 45682 78364
rect 45881 74397 45999 78331
rect 46270 74364 46330 78364
rect 46530 74364 46602 78364
rect 46801 74397 46919 78331
rect 47190 74364 47250 78364
rect 47450 74364 47522 78364
rect 47721 74397 47839 78331
rect 48110 74364 48170 78364
rect 48370 74364 48442 78364
rect 48641 74397 48759 78331
rect 49030 74364 49090 78364
rect 49290 74364 49362 78364
rect 49561 74397 49679 78331
rect 49950 74364 50010 78364
rect 50210 74364 50282 78364
rect 50481 74397 50599 78331
rect 50870 74364 50930 78364
rect 63201 77804 63202 77828
rect 63282 77804 63283 77828
rect 64037 77804 64038 77828
rect 64118 77804 64119 77828
rect 64873 77804 64874 77828
rect 64954 77804 64955 77828
rect 65709 77804 65710 77828
rect 65790 77804 65791 77828
rect 66545 77804 66546 77828
rect 66626 77804 66627 77828
rect 67381 77804 67382 77828
rect 67462 77804 67463 77828
rect 68217 77804 68218 77828
rect 68298 77804 68299 77828
rect 69053 77804 69054 77828
rect 69134 77804 69135 77828
rect 69889 77804 69890 77828
rect 69970 77804 69971 77828
rect 70725 77804 70726 77828
rect 70806 77804 70807 77828
rect 71561 77804 71562 77828
rect 71642 77804 71643 77828
rect 72397 77804 72398 77828
rect 72478 77804 72479 77828
rect 73233 77804 73234 77828
rect 73314 77804 73315 77828
rect 63225 77780 63259 77792
rect 64061 77780 64095 77792
rect 64897 77780 64931 77792
rect 65733 77780 65767 77792
rect 66569 77780 66603 77792
rect 67405 77780 67439 77792
rect 68241 77780 68275 77792
rect 69077 77780 69111 77792
rect 69913 77780 69947 77792
rect 70749 77780 70783 77792
rect 71585 77780 71619 77792
rect 72421 77780 72455 77792
rect 73257 77780 73291 77792
rect 82203 77610 82204 77634
rect 82284 77610 82285 77634
rect 83039 77610 83040 77634
rect 83120 77610 83121 77634
rect 83875 77610 83876 77634
rect 83956 77610 83957 77634
rect 84711 77610 84712 77634
rect 84792 77610 84793 77634
rect 85547 77610 85548 77634
rect 85628 77610 85629 77634
rect 86383 77610 86384 77634
rect 86464 77610 86465 77634
rect 87219 77610 87220 77634
rect 87300 77610 87301 77634
rect 88055 77610 88056 77634
rect 88136 77610 88137 77634
rect 88891 77610 88892 77634
rect 88972 77610 88973 77634
rect 89727 77610 89728 77634
rect 89808 77610 89809 77634
rect 90563 77610 90564 77634
rect 90644 77610 90645 77634
rect 91399 77610 91400 77634
rect 91480 77610 91481 77634
rect 92235 77610 92236 77634
rect 92316 77610 92317 77634
rect 82227 77586 82261 77598
rect 83063 77586 83097 77598
rect 83899 77586 83933 77598
rect 84735 77586 84769 77598
rect 85571 77586 85605 77598
rect 86407 77586 86441 77598
rect 87243 77586 87277 77598
rect 88079 77586 88113 77598
rect 88915 77586 88949 77598
rect 89751 77586 89785 77598
rect 90587 77586 90621 77598
rect 91423 77586 91457 77598
rect 92259 77586 92293 77598
rect 103638 76996 103710 80996
rect 103909 77029 104027 80963
rect 104298 76996 104358 80996
rect 104558 76996 104630 80996
rect 104829 77029 104947 80963
rect 105218 76996 105278 80996
rect 105478 76996 105550 80996
rect 105749 77029 105867 80963
rect 106138 76996 106198 80996
rect 106398 76996 106470 80996
rect 106669 77029 106787 80963
rect 107058 76996 107118 80996
rect 107318 76996 107390 80996
rect 107589 77029 107707 80963
rect 107978 76996 108038 80996
rect 108238 76996 108310 80996
rect 108509 77029 108627 80963
rect 108898 76996 108958 80996
rect 109158 76996 109230 80996
rect 109429 77029 109547 80963
rect 109818 76996 109878 80996
rect 110078 76996 110150 80996
rect 110349 77029 110467 80963
rect 110738 76996 110798 80996
rect 110998 76996 111070 80996
rect 111269 77029 111387 80963
rect 111658 76996 111718 80996
rect 111918 76996 111990 80996
rect 112189 77029 112307 80963
rect 112578 76996 112638 80996
rect 112838 76996 112910 80996
rect 113109 77029 113227 80963
rect 113498 76996 113558 80996
rect 63201 75804 63202 75828
rect 63282 75804 63283 75828
rect 64037 75804 64038 75828
rect 64118 75804 64119 75828
rect 64873 75804 64874 75828
rect 64954 75804 64955 75828
rect 65709 75804 65710 75828
rect 65790 75804 65791 75828
rect 66545 75804 66546 75828
rect 66626 75804 66627 75828
rect 67381 75804 67382 75828
rect 67462 75804 67463 75828
rect 68217 75804 68218 75828
rect 68298 75804 68299 75828
rect 69053 75804 69054 75828
rect 69134 75804 69135 75828
rect 69889 75804 69890 75828
rect 69970 75804 69971 75828
rect 70725 75804 70726 75828
rect 70806 75804 70807 75828
rect 71561 75804 71562 75828
rect 71642 75804 71643 75828
rect 72397 75804 72398 75828
rect 72478 75804 72479 75828
rect 73233 75804 73234 75828
rect 73314 75804 73315 75828
rect 63225 75780 63259 75792
rect 64061 75780 64095 75792
rect 64897 75780 64931 75792
rect 65733 75780 65767 75792
rect 66569 75780 66603 75792
rect 67405 75780 67439 75792
rect 68241 75780 68275 75792
rect 69077 75780 69111 75792
rect 69913 75780 69947 75792
rect 70749 75780 70783 75792
rect 71585 75780 71619 75792
rect 72421 75780 72455 75792
rect 73257 75780 73291 75792
rect 82203 75610 82204 75634
rect 82284 75610 82285 75634
rect 83039 75610 83040 75634
rect 83120 75610 83121 75634
rect 83875 75610 83876 75634
rect 83956 75610 83957 75634
rect 84711 75610 84712 75634
rect 84792 75610 84793 75634
rect 85547 75610 85548 75634
rect 85628 75610 85629 75634
rect 86383 75610 86384 75634
rect 86464 75610 86465 75634
rect 87219 75610 87220 75634
rect 87300 75610 87301 75634
rect 88055 75610 88056 75634
rect 88136 75610 88137 75634
rect 88891 75610 88892 75634
rect 88972 75610 88973 75634
rect 89727 75610 89728 75634
rect 89808 75610 89809 75634
rect 90563 75610 90564 75634
rect 90644 75610 90645 75634
rect 91399 75610 91400 75634
rect 91480 75610 91481 75634
rect 92235 75610 92236 75634
rect 92316 75610 92317 75634
rect 82227 75586 82261 75598
rect 83063 75586 83097 75598
rect 83899 75586 83933 75598
rect 84735 75586 84769 75598
rect 85571 75586 85605 75598
rect 86407 75586 86441 75598
rect 87243 75586 87277 75598
rect 88079 75586 88113 75598
rect 88915 75586 88949 75598
rect 89751 75586 89785 75598
rect 90587 75586 90621 75598
rect 91423 75586 91457 75598
rect 92259 75586 92293 75598
rect 63201 73804 63202 73828
rect 63282 73804 63283 73828
rect 64037 73804 64038 73828
rect 64118 73804 64119 73828
rect 64873 73804 64874 73828
rect 64954 73804 64955 73828
rect 65709 73804 65710 73828
rect 65790 73804 65791 73828
rect 66545 73804 66546 73828
rect 66626 73804 66627 73828
rect 67381 73804 67382 73828
rect 67462 73804 67463 73828
rect 68217 73804 68218 73828
rect 68298 73804 68299 73828
rect 69053 73804 69054 73828
rect 69134 73804 69135 73828
rect 69889 73804 69890 73828
rect 69970 73804 69971 73828
rect 70725 73804 70726 73828
rect 70806 73804 70807 73828
rect 71561 73804 71562 73828
rect 71642 73804 71643 73828
rect 72397 73804 72398 73828
rect 72478 73804 72479 73828
rect 73233 73804 73234 73828
rect 73314 73804 73315 73828
rect 63225 73780 63259 73792
rect 64061 73780 64095 73792
rect 64897 73780 64931 73792
rect 65733 73780 65767 73792
rect 66569 73780 66603 73792
rect 67405 73780 67439 73792
rect 68241 73780 68275 73792
rect 69077 73780 69111 73792
rect 69913 73780 69947 73792
rect 70749 73780 70783 73792
rect 71585 73780 71619 73792
rect 72421 73780 72455 73792
rect 73257 73780 73291 73792
rect 4377 73550 4378 73574
rect 4458 73550 4459 73574
rect 5213 73550 5214 73574
rect 5294 73550 5295 73574
rect 6049 73550 6050 73574
rect 6130 73550 6131 73574
rect 6885 73550 6886 73574
rect 6966 73550 6967 73574
rect 7721 73550 7722 73574
rect 7802 73550 7803 73574
rect 8557 73550 8558 73574
rect 8638 73550 8639 73574
rect 9393 73550 9394 73574
rect 9474 73550 9475 73574
rect 10229 73550 10230 73574
rect 10310 73550 10311 73574
rect 11065 73550 11066 73574
rect 11146 73550 11147 73574
rect 11901 73550 11902 73574
rect 11982 73550 11983 73574
rect 12737 73550 12738 73574
rect 12818 73550 12819 73574
rect 4401 73526 4435 73538
rect 5237 73526 5271 73538
rect 6073 73526 6107 73538
rect 6909 73526 6943 73538
rect 7745 73526 7779 73538
rect 8581 73526 8615 73538
rect 9417 73526 9451 73538
rect 10253 73526 10287 73538
rect 11089 73526 11123 73538
rect 11925 73526 11959 73538
rect 12761 73526 12795 73538
rect 4377 71929 4378 71953
rect 4458 71929 4459 71953
rect 5213 71929 5214 71953
rect 5294 71929 5295 71953
rect 6049 71929 6050 71953
rect 6130 71929 6131 71953
rect 6885 71929 6886 71953
rect 6966 71929 6967 71953
rect 7721 71929 7722 71953
rect 7802 71929 7803 71953
rect 8557 71929 8558 71953
rect 8638 71929 8639 71953
rect 9393 71929 9394 71953
rect 9474 71929 9475 71953
rect 10229 71929 10230 71953
rect 10310 71929 10311 71953
rect 11065 71929 11066 71953
rect 11146 71929 11147 71953
rect 11901 71929 11902 71953
rect 11982 71929 11983 71953
rect 12737 71929 12738 71953
rect 12818 71929 12819 71953
rect 4401 71905 4435 71917
rect 5237 71905 5271 71917
rect 6073 71905 6107 71917
rect 6909 71905 6943 71917
rect 7745 71905 7779 71917
rect 8581 71905 8615 71917
rect 9417 71905 9451 71917
rect 10253 71905 10287 71917
rect 11089 71905 11123 71917
rect 11925 71905 11959 71917
rect 12761 71905 12795 71917
rect 23072 69570 23144 73570
rect 23343 69603 23461 73537
rect 23732 69570 23792 73570
rect 23992 69570 24064 73570
rect 24263 69603 24381 73537
rect 24652 69570 24712 73570
rect 24912 69570 24984 73570
rect 25183 69603 25301 73537
rect 25572 69570 25632 73570
rect 25832 69570 25904 73570
rect 26103 69603 26221 73537
rect 26492 69570 26552 73570
rect 26752 69570 26824 73570
rect 27023 69603 27141 73537
rect 27412 69570 27472 73570
rect 27672 69570 27744 73570
rect 27943 69603 28061 73537
rect 28332 69570 28392 73570
rect 28592 69570 28664 73570
rect 28863 69603 28981 73537
rect 29252 69570 29312 73570
rect 29512 69570 29584 73570
rect 29783 69603 29901 73537
rect 30172 69570 30232 73570
rect 30432 69570 30504 73570
rect 30703 69603 30821 73537
rect 31092 69570 31152 73570
rect 42850 69764 42922 73764
rect 43121 69797 43239 73731
rect 43510 69764 43570 73764
rect 43770 69764 43842 73764
rect 44041 69797 44159 73731
rect 44430 69764 44490 73764
rect 44690 69764 44762 73764
rect 44961 69797 45079 73731
rect 45350 69764 45410 73764
rect 45610 69764 45682 73764
rect 45881 69797 45999 73731
rect 46270 69764 46330 73764
rect 46530 69764 46602 73764
rect 46801 69797 46919 73731
rect 47190 69764 47250 73764
rect 47450 69764 47522 73764
rect 47721 69797 47839 73731
rect 48110 69764 48170 73764
rect 48370 69764 48442 73764
rect 48641 69797 48759 73731
rect 49030 69764 49090 73764
rect 49290 69764 49362 73764
rect 49561 69797 49679 73731
rect 49950 69764 50010 73764
rect 50210 69764 50282 73764
rect 50481 69797 50599 73731
rect 50870 69764 50930 73764
rect 82203 73610 82204 73634
rect 82284 73610 82285 73634
rect 83039 73610 83040 73634
rect 83120 73610 83121 73634
rect 83875 73610 83876 73634
rect 83956 73610 83957 73634
rect 84711 73610 84712 73634
rect 84792 73610 84793 73634
rect 85547 73610 85548 73634
rect 85628 73610 85629 73634
rect 86383 73610 86384 73634
rect 86464 73610 86465 73634
rect 87219 73610 87220 73634
rect 87300 73610 87301 73634
rect 88055 73610 88056 73634
rect 88136 73610 88137 73634
rect 88891 73610 88892 73634
rect 88972 73610 88973 73634
rect 89727 73610 89728 73634
rect 89808 73610 89809 73634
rect 90563 73610 90564 73634
rect 90644 73610 90645 73634
rect 91399 73610 91400 73634
rect 91480 73610 91481 73634
rect 92235 73610 92236 73634
rect 92316 73610 92317 73634
rect 82227 73586 82261 73598
rect 83063 73586 83097 73598
rect 83899 73586 83933 73598
rect 84735 73586 84769 73598
rect 85571 73586 85605 73598
rect 86407 73586 86441 73598
rect 87243 73586 87277 73598
rect 88079 73586 88113 73598
rect 88915 73586 88949 73598
rect 89751 73586 89785 73598
rect 90587 73586 90621 73598
rect 91423 73586 91457 73598
rect 92259 73586 92293 73598
rect 103638 72396 103710 76396
rect 103909 72429 104027 76363
rect 104298 72396 104358 76396
rect 104558 72396 104630 76396
rect 104829 72429 104947 76363
rect 105218 72396 105278 76396
rect 105478 72396 105550 76396
rect 105749 72429 105867 76363
rect 106138 72396 106198 76396
rect 106398 72396 106470 76396
rect 106669 72429 106787 76363
rect 107058 72396 107118 76396
rect 107318 72396 107390 76396
rect 107589 72429 107707 76363
rect 107978 72396 108038 76396
rect 108238 72396 108310 76396
rect 108509 72429 108627 76363
rect 108898 72396 108958 76396
rect 109158 72396 109230 76396
rect 109429 72429 109547 76363
rect 109818 72396 109878 76396
rect 110078 72396 110150 76396
rect 110349 72429 110467 76363
rect 110738 72396 110798 76396
rect 110998 72396 111070 76396
rect 111269 72429 111387 76363
rect 111658 72396 111718 76396
rect 111918 72396 111990 76396
rect 112189 72429 112307 76363
rect 112578 72396 112638 76396
rect 112838 72396 112910 76396
rect 113109 72429 113227 76363
rect 113498 72396 113558 76396
rect 64873 71804 64874 71828
rect 64954 71804 64955 71828
rect 65709 71804 65710 71828
rect 65790 71804 65791 71828
rect 66545 71804 66546 71828
rect 66626 71804 66627 71828
rect 67381 71804 67382 71828
rect 67462 71804 67463 71828
rect 68217 71804 68218 71828
rect 68298 71804 68299 71828
rect 69053 71804 69054 71828
rect 69134 71804 69135 71828
rect 69889 71804 69890 71828
rect 69970 71804 69971 71828
rect 70725 71804 70726 71828
rect 70806 71804 70807 71828
rect 71561 71804 71562 71828
rect 71642 71804 71643 71828
rect 72397 71804 72398 71828
rect 72478 71804 72479 71828
rect 73233 71804 73234 71828
rect 73314 71804 73315 71828
rect 64897 71780 64931 71792
rect 65733 71780 65767 71792
rect 66569 71780 66603 71792
rect 67405 71780 67439 71792
rect 68241 71780 68275 71792
rect 69077 71780 69111 71792
rect 69913 71780 69947 71792
rect 70749 71780 70783 71792
rect 71585 71780 71619 71792
rect 72421 71780 72455 71792
rect 73257 71780 73291 71792
rect 83875 71610 83876 71634
rect 83956 71610 83957 71634
rect 84711 71610 84712 71634
rect 84792 71610 84793 71634
rect 85547 71610 85548 71634
rect 85628 71610 85629 71634
rect 86383 71610 86384 71634
rect 86464 71610 86465 71634
rect 87219 71610 87220 71634
rect 87300 71610 87301 71634
rect 88055 71610 88056 71634
rect 88136 71610 88137 71634
rect 88891 71610 88892 71634
rect 88972 71610 88973 71634
rect 89727 71610 89728 71634
rect 89808 71610 89809 71634
rect 90563 71610 90564 71634
rect 90644 71610 90645 71634
rect 91399 71610 91400 71634
rect 91480 71610 91481 71634
rect 92235 71610 92236 71634
rect 92316 71610 92317 71634
rect 83899 71586 83933 71598
rect 84735 71586 84769 71598
rect 85571 71586 85605 71598
rect 86407 71586 86441 71598
rect 87243 71586 87277 71598
rect 88079 71586 88113 71598
rect 88915 71586 88949 71598
rect 89751 71586 89785 71598
rect 90587 71586 90621 71598
rect 91423 71586 91457 71598
rect 92259 71586 92293 71598
rect 64873 70183 64874 70207
rect 64954 70183 64955 70207
rect 65709 70183 65710 70207
rect 65790 70183 65791 70207
rect 66545 70183 66546 70207
rect 66626 70183 66627 70207
rect 67381 70183 67382 70207
rect 67462 70183 67463 70207
rect 68217 70183 68218 70207
rect 68298 70183 68299 70207
rect 69053 70183 69054 70207
rect 69134 70183 69135 70207
rect 69889 70183 69890 70207
rect 69970 70183 69971 70207
rect 70725 70183 70726 70207
rect 70806 70183 70807 70207
rect 71561 70183 71562 70207
rect 71642 70183 71643 70207
rect 72397 70183 72398 70207
rect 72478 70183 72479 70207
rect 73233 70183 73234 70207
rect 73314 70183 73315 70207
rect 64897 70159 64931 70171
rect 65733 70159 65767 70171
rect 66569 70159 66603 70171
rect 67405 70159 67439 70171
rect 68241 70159 68275 70171
rect 69077 70159 69111 70171
rect 69913 70159 69947 70171
rect 70749 70159 70783 70171
rect 71585 70159 71619 70171
rect 72421 70159 72455 70171
rect 73257 70159 73291 70171
rect 83875 69989 83876 70013
rect 83956 69989 83957 70013
rect 84711 69989 84712 70013
rect 84792 69989 84793 70013
rect 85547 69989 85548 70013
rect 85628 69989 85629 70013
rect 86383 69989 86384 70013
rect 86464 69989 86465 70013
rect 87219 69989 87220 70013
rect 87300 69989 87301 70013
rect 88055 69989 88056 70013
rect 88136 69989 88137 70013
rect 88891 69989 88892 70013
rect 88972 69989 88973 70013
rect 89727 69989 89728 70013
rect 89808 69989 89809 70013
rect 90563 69989 90564 70013
rect 90644 69989 90645 70013
rect 91399 69989 91400 70013
rect 91480 69989 91481 70013
rect 92235 69989 92236 70013
rect 92316 69989 92317 70013
rect 83899 69965 83933 69977
rect 84735 69965 84769 69977
rect 85571 69965 85605 69977
rect 86407 69965 86441 69977
rect 87243 69965 87277 69977
rect 88079 69965 88113 69977
rect 88915 69965 88949 69977
rect 89751 69965 89785 69977
rect 90587 69965 90621 69977
rect 91423 69965 91457 69977
rect 92259 69965 92293 69977
rect 23072 64970 23144 68970
rect 23343 65003 23461 68937
rect 23732 64970 23792 68970
rect 23992 64970 24064 68970
rect 24263 65003 24381 68937
rect 24652 64970 24712 68970
rect 24912 64970 24984 68970
rect 25183 65003 25301 68937
rect 25572 64970 25632 68970
rect 25832 64970 25904 68970
rect 26103 65003 26221 68937
rect 26492 64970 26552 68970
rect 26752 64970 26824 68970
rect 27023 65003 27141 68937
rect 27412 64970 27472 68970
rect 27672 64970 27744 68970
rect 27943 65003 28061 68937
rect 28332 64970 28392 68970
rect 28592 64970 28664 68970
rect 28863 65003 28981 68937
rect 29252 64970 29312 68970
rect 29512 64970 29584 68970
rect 29783 65003 29901 68937
rect 30172 64970 30232 68970
rect 30432 64970 30504 68970
rect 30703 65003 30821 68937
rect 31092 64970 31152 68970
rect 42850 65164 42922 69164
rect 43121 65197 43239 69131
rect 43510 65164 43570 69164
rect 43770 65164 43842 69164
rect 44041 65197 44159 69131
rect 44430 65164 44490 69164
rect 44690 65164 44762 69164
rect 44961 65197 45079 69131
rect 45350 65164 45410 69164
rect 45610 65164 45682 69164
rect 45881 65197 45999 69131
rect 46270 65164 46330 69164
rect 46530 65164 46602 69164
rect 46801 65197 46919 69131
rect 47190 65164 47250 69164
rect 47450 65164 47522 69164
rect 47721 65197 47839 69131
rect 48110 65164 48170 69164
rect 48370 65164 48442 69164
rect 48641 65197 48759 69131
rect 49030 65164 49090 69164
rect 49290 65164 49362 69164
rect 49561 65197 49679 69131
rect 49950 65164 50010 69164
rect 50210 65164 50282 69164
rect 50481 65197 50599 69131
rect 50870 65164 50930 69164
rect 105478 67796 105550 71796
rect 105749 67829 105867 71763
rect 106138 67796 106198 71796
rect 106398 67796 106470 71796
rect 106669 67829 106787 71763
rect 107058 67796 107118 71796
rect 107318 67796 107390 71796
rect 107589 67829 107707 71763
rect 107978 67796 108038 71796
rect 108238 67796 108310 71796
rect 108509 67829 108627 71763
rect 108898 67796 108958 71796
rect 109158 67796 109230 71796
rect 109429 67829 109547 71763
rect 109818 67796 109878 71796
rect 110078 67796 110150 71796
rect 110349 67829 110467 71763
rect 110738 67796 110798 71796
rect 110998 67796 111070 71796
rect 111269 67829 111387 71763
rect 111658 67796 111718 71796
rect 111918 67796 111990 71796
rect 112189 67829 112307 71763
rect 112578 67796 112638 71796
rect 112838 67796 112910 71796
rect 113109 67829 113227 71763
rect 113498 67796 113558 71796
rect 23072 60370 23144 64370
rect 23343 60403 23461 64337
rect 23732 60370 23792 64370
rect 23992 60370 24064 64370
rect 24263 60403 24381 64337
rect 24652 60370 24712 64370
rect 24912 60370 24984 64370
rect 25183 60403 25301 64337
rect 25572 60370 25632 64370
rect 25832 60370 25904 64370
rect 26103 60403 26221 64337
rect 26492 60370 26552 64370
rect 26752 60370 26824 64370
rect 27023 60403 27141 64337
rect 27412 60370 27472 64370
rect 27672 60370 27744 64370
rect 27943 60403 28061 64337
rect 28332 60370 28392 64370
rect 28592 60370 28664 64370
rect 28863 60403 28981 64337
rect 29252 60370 29312 64370
rect 29512 60370 29584 64370
rect 29783 60403 29901 64337
rect 30172 60370 30232 64370
rect 30432 60370 30504 64370
rect 30703 60403 30821 64337
rect 31092 60370 31152 64370
rect 42850 60564 42922 64564
rect 43121 60597 43239 64531
rect 43510 60564 43570 64564
rect 43770 60564 43842 64564
rect 44041 60597 44159 64531
rect 44430 60564 44490 64564
rect 44690 60564 44762 64564
rect 44961 60597 45079 64531
rect 45350 60564 45410 64564
rect 45610 60564 45682 64564
rect 45881 60597 45999 64531
rect 46270 60564 46330 64564
rect 46530 60564 46602 64564
rect 46801 60597 46919 64531
rect 47190 60564 47250 64564
rect 47450 60564 47522 64564
rect 47721 60597 47839 64531
rect 48110 60564 48170 64564
rect 48370 60564 48442 64564
rect 48641 60597 48759 64531
rect 49030 60564 49090 64564
rect 49290 60564 49362 64564
rect 49561 60597 49679 64531
rect 49950 60564 50010 64564
rect 50210 60564 50282 64564
rect 50481 60597 50599 64531
rect 50870 60564 50930 64564
rect 105478 63196 105550 67196
rect 105749 63229 105867 67163
rect 106138 63196 106198 67196
rect 106398 63196 106470 67196
rect 106669 63229 106787 67163
rect 107058 63196 107118 67196
rect 107318 63196 107390 67196
rect 107589 63229 107707 67163
rect 107978 63196 108038 67196
rect 108238 63196 108310 67196
rect 108509 63229 108627 67163
rect 108898 63196 108958 67196
rect 109158 63196 109230 67196
rect 109429 63229 109547 67163
rect 109818 63196 109878 67196
rect 110078 63196 110150 67196
rect 110349 63229 110467 67163
rect 110738 63196 110798 67196
rect 110998 63196 111070 67196
rect 111269 63229 111387 67163
rect 111658 63196 111718 67196
rect 111918 63196 111990 67196
rect 112189 63229 112307 67163
rect 112578 63196 112638 67196
rect 112838 63196 112910 67196
rect 113109 63229 113227 67163
rect 113498 63196 113558 67196
rect 2211 59550 2212 59574
rect 2292 59550 2293 59574
rect 2765 59550 2766 59574
rect 2846 59550 2847 59574
rect 3319 59550 3320 59574
rect 3400 59550 3401 59574
rect 3873 59550 3874 59574
rect 3954 59550 3955 59574
rect 4427 59550 4428 59574
rect 4508 59550 4509 59574
rect 4981 59550 4982 59574
rect 5062 59550 5063 59574
rect 5535 59550 5536 59574
rect 5616 59550 5617 59574
rect 6089 59550 6090 59574
rect 6170 59550 6171 59574
rect 6643 59550 6644 59574
rect 6724 59550 6725 59574
rect 7197 59550 7198 59574
rect 7278 59550 7279 59574
rect 7751 59550 7752 59574
rect 7832 59550 7833 59574
rect 8305 59550 8306 59574
rect 8386 59550 8387 59574
rect 8859 59550 8860 59574
rect 8940 59550 8941 59574
rect 9413 59550 9414 59574
rect 9494 59550 9495 59574
rect 9967 59550 9968 59574
rect 10048 59550 10049 59574
rect 10521 59550 10522 59574
rect 10602 59550 10603 59574
rect 11075 59550 11076 59574
rect 11156 59550 11157 59574
rect 11629 59550 11630 59574
rect 11710 59550 11711 59574
rect 12183 59550 12184 59574
rect 12264 59550 12265 59574
rect 12737 59550 12738 59574
rect 12818 59550 12819 59574
rect 2235 59526 2269 59538
rect 2789 59526 2823 59538
rect 3343 59526 3377 59538
rect 3897 59526 3931 59538
rect 4451 59526 4485 59538
rect 5005 59526 5039 59538
rect 5559 59526 5593 59538
rect 6113 59526 6147 59538
rect 6667 59526 6701 59538
rect 7221 59526 7255 59538
rect 7775 59526 7809 59538
rect 8329 59526 8363 59538
rect 8883 59526 8917 59538
rect 9437 59526 9471 59538
rect 9991 59526 10025 59538
rect 10545 59526 10579 59538
rect 11099 59526 11133 59538
rect 11653 59526 11687 59538
rect 12207 59526 12241 59538
rect 12761 59526 12795 59538
rect 2211 57550 2212 57574
rect 2292 57550 2293 57574
rect 2765 57550 2766 57574
rect 2846 57550 2847 57574
rect 3319 57550 3320 57574
rect 3400 57550 3401 57574
rect 3873 57550 3874 57574
rect 3954 57550 3955 57574
rect 4427 57550 4428 57574
rect 4508 57550 4509 57574
rect 4981 57550 4982 57574
rect 5062 57550 5063 57574
rect 5535 57550 5536 57574
rect 5616 57550 5617 57574
rect 6089 57550 6090 57574
rect 6170 57550 6171 57574
rect 6643 57550 6644 57574
rect 6724 57550 6725 57574
rect 7197 57550 7198 57574
rect 7278 57550 7279 57574
rect 7751 57550 7752 57574
rect 7832 57550 7833 57574
rect 8305 57550 8306 57574
rect 8386 57550 8387 57574
rect 8859 57550 8860 57574
rect 8940 57550 8941 57574
rect 9413 57550 9414 57574
rect 9494 57550 9495 57574
rect 9967 57550 9968 57574
rect 10048 57550 10049 57574
rect 10521 57550 10522 57574
rect 10602 57550 10603 57574
rect 11075 57550 11076 57574
rect 11156 57550 11157 57574
rect 11629 57550 11630 57574
rect 11710 57550 11711 57574
rect 12183 57550 12184 57574
rect 12264 57550 12265 57574
rect 12737 57550 12738 57574
rect 12818 57550 12819 57574
rect 2235 57526 2269 57538
rect 2789 57526 2823 57538
rect 3343 57526 3377 57538
rect 3897 57526 3931 57538
rect 4451 57526 4485 57538
rect 5005 57526 5039 57538
rect 5559 57526 5593 57538
rect 6113 57526 6147 57538
rect 6667 57526 6701 57538
rect 7221 57526 7255 57538
rect 7775 57526 7809 57538
rect 8329 57526 8363 57538
rect 8883 57526 8917 57538
rect 9437 57526 9471 57538
rect 9991 57526 10025 57538
rect 10545 57526 10579 57538
rect 11099 57526 11133 57538
rect 11653 57526 11687 57538
rect 12207 57526 12241 57538
rect 12761 57526 12795 57538
rect 21232 55770 21304 59770
rect 21503 55803 21621 59737
rect 21892 55770 21952 59770
rect 22152 55770 22224 59770
rect 22423 55803 22541 59737
rect 22812 55770 22872 59770
rect 23072 55770 23144 59770
rect 23343 55803 23461 59737
rect 23732 55770 23792 59770
rect 23992 55770 24064 59770
rect 24263 55803 24381 59737
rect 24652 55770 24712 59770
rect 24912 55770 24984 59770
rect 25183 55803 25301 59737
rect 25572 55770 25632 59770
rect 25832 55770 25904 59770
rect 26103 55803 26221 59737
rect 26492 55770 26552 59770
rect 26752 55770 26824 59770
rect 27023 55803 27141 59737
rect 27412 55770 27472 59770
rect 27672 55770 27744 59770
rect 27943 55803 28061 59737
rect 28332 55770 28392 59770
rect 28592 55770 28664 59770
rect 28863 55803 28981 59737
rect 29252 55770 29312 59770
rect 29512 55770 29584 59770
rect 29783 55803 29901 59737
rect 30172 55770 30232 59770
rect 30432 55770 30504 59770
rect 30703 55803 30821 59737
rect 31092 55770 31152 59770
rect 41010 55964 41082 59964
rect 41281 55997 41399 59931
rect 41670 55964 41730 59964
rect 41930 55964 42002 59964
rect 42201 55997 42319 59931
rect 42590 55964 42650 59964
rect 42850 55964 42922 59964
rect 43121 55997 43239 59931
rect 43510 55964 43570 59964
rect 43770 55964 43842 59964
rect 44041 55997 44159 59931
rect 44430 55964 44490 59964
rect 44690 55964 44762 59964
rect 44961 55997 45079 59931
rect 45350 55964 45410 59964
rect 45610 55964 45682 59964
rect 45881 55997 45999 59931
rect 46270 55964 46330 59964
rect 46530 55964 46602 59964
rect 46801 55997 46919 59931
rect 47190 55964 47250 59964
rect 47450 55964 47522 59964
rect 47721 55997 47839 59931
rect 48110 55964 48170 59964
rect 48370 55964 48442 59964
rect 48641 55997 48759 59931
rect 49030 55964 49090 59964
rect 49290 55964 49362 59964
rect 49561 55997 49679 59931
rect 49950 55964 50010 59964
rect 50210 55964 50282 59964
rect 50481 55997 50599 59931
rect 50870 55964 50930 59964
rect 105478 58596 105550 62596
rect 105749 58629 105867 62563
rect 106138 58596 106198 62596
rect 106398 58596 106470 62596
rect 106669 58629 106787 62563
rect 107058 58596 107118 62596
rect 107318 58596 107390 62596
rect 107589 58629 107707 62563
rect 107978 58596 108038 62596
rect 108238 58596 108310 62596
rect 108509 58629 108627 62563
rect 108898 58596 108958 62596
rect 109158 58596 109230 62596
rect 109429 58629 109547 62563
rect 109818 58596 109878 62596
rect 110078 58596 110150 62596
rect 110349 58629 110467 62563
rect 110738 58596 110798 62596
rect 110998 58596 111070 62596
rect 111269 58629 111387 62563
rect 111658 58596 111718 62596
rect 111918 58596 111990 62596
rect 112189 58629 112307 62563
rect 112578 58596 112638 62596
rect 112838 58596 112910 62596
rect 113109 58629 113227 62563
rect 113498 58596 113558 62596
rect 62707 57804 62708 57828
rect 62788 57804 62789 57828
rect 63261 57804 63262 57828
rect 63342 57804 63343 57828
rect 63815 57804 63816 57828
rect 63896 57804 63897 57828
rect 64369 57804 64370 57828
rect 64450 57804 64451 57828
rect 64923 57804 64924 57828
rect 65004 57804 65005 57828
rect 65477 57804 65478 57828
rect 65558 57804 65559 57828
rect 66031 57804 66032 57828
rect 66112 57804 66113 57828
rect 66585 57804 66586 57828
rect 66666 57804 66667 57828
rect 67139 57804 67140 57828
rect 67220 57804 67221 57828
rect 67693 57804 67694 57828
rect 67774 57804 67775 57828
rect 68247 57804 68248 57828
rect 68328 57804 68329 57828
rect 68801 57804 68802 57828
rect 68882 57804 68883 57828
rect 69355 57804 69356 57828
rect 69436 57804 69437 57828
rect 69909 57804 69910 57828
rect 69990 57804 69991 57828
rect 70463 57804 70464 57828
rect 70544 57804 70545 57828
rect 71017 57804 71018 57828
rect 71098 57804 71099 57828
rect 71571 57804 71572 57828
rect 71652 57804 71653 57828
rect 72125 57804 72126 57828
rect 72206 57804 72207 57828
rect 72679 57804 72680 57828
rect 72760 57804 72761 57828
rect 73233 57804 73234 57828
rect 73314 57804 73315 57828
rect 62731 57780 62765 57792
rect 63285 57780 63319 57792
rect 63839 57780 63873 57792
rect 64393 57780 64427 57792
rect 64947 57780 64981 57792
rect 65501 57780 65535 57792
rect 66055 57780 66089 57792
rect 66609 57780 66643 57792
rect 67163 57780 67197 57792
rect 67717 57780 67751 57792
rect 68271 57780 68305 57792
rect 68825 57780 68859 57792
rect 69379 57780 69413 57792
rect 69933 57780 69967 57792
rect 70487 57780 70521 57792
rect 71041 57780 71075 57792
rect 71595 57780 71629 57792
rect 72149 57780 72183 57792
rect 72703 57780 72737 57792
rect 73257 57780 73291 57792
rect 81709 57610 81710 57634
rect 81790 57610 81791 57634
rect 82263 57610 82264 57634
rect 82344 57610 82345 57634
rect 82817 57610 82818 57634
rect 82898 57610 82899 57634
rect 83371 57610 83372 57634
rect 83452 57610 83453 57634
rect 83925 57610 83926 57634
rect 84006 57610 84007 57634
rect 84479 57610 84480 57634
rect 84560 57610 84561 57634
rect 85033 57610 85034 57634
rect 85114 57610 85115 57634
rect 85587 57610 85588 57634
rect 85668 57610 85669 57634
rect 86141 57610 86142 57634
rect 86222 57610 86223 57634
rect 86695 57610 86696 57634
rect 86776 57610 86777 57634
rect 87249 57610 87250 57634
rect 87330 57610 87331 57634
rect 87803 57610 87804 57634
rect 87884 57610 87885 57634
rect 88357 57610 88358 57634
rect 88438 57610 88439 57634
rect 88911 57610 88912 57634
rect 88992 57610 88993 57634
rect 89465 57610 89466 57634
rect 89546 57610 89547 57634
rect 90019 57610 90020 57634
rect 90100 57610 90101 57634
rect 90573 57610 90574 57634
rect 90654 57610 90655 57634
rect 91127 57610 91128 57634
rect 91208 57610 91209 57634
rect 91681 57610 91682 57634
rect 91762 57610 91763 57634
rect 92235 57610 92236 57634
rect 92316 57610 92317 57634
rect 81733 57586 81767 57598
rect 82287 57586 82321 57598
rect 82841 57586 82875 57598
rect 83395 57586 83429 57598
rect 83949 57586 83983 57598
rect 84503 57586 84537 57598
rect 85057 57586 85091 57598
rect 85611 57586 85645 57598
rect 86165 57586 86199 57598
rect 86719 57586 86753 57598
rect 87273 57586 87307 57598
rect 87827 57586 87861 57598
rect 88381 57586 88415 57598
rect 88935 57586 88969 57598
rect 89489 57586 89523 57598
rect 90043 57586 90077 57598
rect 90597 57586 90631 57598
rect 91151 57586 91185 57598
rect 91705 57586 91739 57598
rect 92259 57586 92293 57598
rect 62707 55804 62708 55828
rect 62788 55804 62789 55828
rect 63261 55804 63262 55828
rect 63342 55804 63343 55828
rect 63815 55804 63816 55828
rect 63896 55804 63897 55828
rect 64369 55804 64370 55828
rect 64450 55804 64451 55828
rect 64923 55804 64924 55828
rect 65004 55804 65005 55828
rect 65477 55804 65478 55828
rect 65558 55804 65559 55828
rect 66031 55804 66032 55828
rect 66112 55804 66113 55828
rect 66585 55804 66586 55828
rect 66666 55804 66667 55828
rect 67139 55804 67140 55828
rect 67220 55804 67221 55828
rect 67693 55804 67694 55828
rect 67774 55804 67775 55828
rect 68247 55804 68248 55828
rect 68328 55804 68329 55828
rect 68801 55804 68802 55828
rect 68882 55804 68883 55828
rect 69355 55804 69356 55828
rect 69436 55804 69437 55828
rect 69909 55804 69910 55828
rect 69990 55804 69991 55828
rect 70463 55804 70464 55828
rect 70544 55804 70545 55828
rect 71017 55804 71018 55828
rect 71098 55804 71099 55828
rect 71571 55804 71572 55828
rect 71652 55804 71653 55828
rect 72125 55804 72126 55828
rect 72206 55804 72207 55828
rect 72679 55804 72680 55828
rect 72760 55804 72761 55828
rect 73233 55804 73234 55828
rect 73314 55804 73315 55828
rect 62731 55780 62765 55792
rect 63285 55780 63319 55792
rect 63839 55780 63873 55792
rect 64393 55780 64427 55792
rect 64947 55780 64981 55792
rect 65501 55780 65535 55792
rect 66055 55780 66089 55792
rect 66609 55780 66643 55792
rect 67163 55780 67197 55792
rect 67717 55780 67751 55792
rect 68271 55780 68305 55792
rect 68825 55780 68859 55792
rect 69379 55780 69413 55792
rect 69933 55780 69967 55792
rect 70487 55780 70521 55792
rect 71041 55780 71075 55792
rect 71595 55780 71629 55792
rect 72149 55780 72183 55792
rect 72703 55780 72737 55792
rect 73257 55780 73291 55792
rect 81709 55610 81710 55634
rect 81790 55610 81791 55634
rect 82263 55610 82264 55634
rect 82344 55610 82345 55634
rect 82817 55610 82818 55634
rect 82898 55610 82899 55634
rect 83371 55610 83372 55634
rect 83452 55610 83453 55634
rect 83925 55610 83926 55634
rect 84006 55610 84007 55634
rect 84479 55610 84480 55634
rect 84560 55610 84561 55634
rect 85033 55610 85034 55634
rect 85114 55610 85115 55634
rect 85587 55610 85588 55634
rect 85668 55610 85669 55634
rect 86141 55610 86142 55634
rect 86222 55610 86223 55634
rect 86695 55610 86696 55634
rect 86776 55610 86777 55634
rect 87249 55610 87250 55634
rect 87330 55610 87331 55634
rect 87803 55610 87804 55634
rect 87884 55610 87885 55634
rect 88357 55610 88358 55634
rect 88438 55610 88439 55634
rect 88911 55610 88912 55634
rect 88992 55610 88993 55634
rect 89465 55610 89466 55634
rect 89546 55610 89547 55634
rect 90019 55610 90020 55634
rect 90100 55610 90101 55634
rect 90573 55610 90574 55634
rect 90654 55610 90655 55634
rect 91127 55610 91128 55634
rect 91208 55610 91209 55634
rect 91681 55610 91682 55634
rect 91762 55610 91763 55634
rect 92235 55610 92236 55634
rect 92316 55610 92317 55634
rect 81733 55586 81767 55598
rect 82287 55586 82321 55598
rect 82841 55586 82875 55598
rect 83395 55586 83429 55598
rect 83949 55586 83983 55598
rect 84503 55586 84537 55598
rect 85057 55586 85091 55598
rect 85611 55586 85645 55598
rect 86165 55586 86199 55598
rect 86719 55586 86753 55598
rect 87273 55586 87307 55598
rect 87827 55586 87861 55598
rect 88381 55586 88415 55598
rect 88935 55586 88969 55598
rect 89489 55586 89523 55598
rect 90043 55586 90077 55598
rect 90597 55586 90631 55598
rect 91151 55586 91185 55598
rect 91705 55586 91739 55598
rect 92259 55586 92293 55598
rect 2211 55550 2212 55574
rect 2292 55550 2293 55574
rect 2765 55550 2766 55574
rect 2846 55550 2847 55574
rect 3319 55550 3320 55574
rect 3400 55550 3401 55574
rect 3873 55550 3874 55574
rect 3954 55550 3955 55574
rect 4427 55550 4428 55574
rect 4508 55550 4509 55574
rect 4981 55550 4982 55574
rect 5062 55550 5063 55574
rect 5535 55550 5536 55574
rect 5616 55550 5617 55574
rect 6089 55550 6090 55574
rect 6170 55550 6171 55574
rect 6643 55550 6644 55574
rect 6724 55550 6725 55574
rect 7197 55550 7198 55574
rect 7278 55550 7279 55574
rect 7751 55550 7752 55574
rect 7832 55550 7833 55574
rect 8305 55550 8306 55574
rect 8386 55550 8387 55574
rect 8859 55550 8860 55574
rect 8940 55550 8941 55574
rect 9413 55550 9414 55574
rect 9494 55550 9495 55574
rect 9967 55550 9968 55574
rect 10048 55550 10049 55574
rect 10521 55550 10522 55574
rect 10602 55550 10603 55574
rect 11075 55550 11076 55574
rect 11156 55550 11157 55574
rect 11629 55550 11630 55574
rect 11710 55550 11711 55574
rect 12183 55550 12184 55574
rect 12264 55550 12265 55574
rect 12737 55550 12738 55574
rect 12818 55550 12819 55574
rect 2235 55526 2269 55538
rect 2789 55526 2823 55538
rect 3343 55526 3377 55538
rect 3897 55526 3931 55538
rect 4451 55526 4485 55538
rect 5005 55526 5039 55538
rect 5559 55526 5593 55538
rect 6113 55526 6147 55538
rect 6667 55526 6701 55538
rect 7221 55526 7255 55538
rect 7775 55526 7809 55538
rect 8329 55526 8363 55538
rect 8883 55526 8917 55538
rect 9437 55526 9471 55538
rect 9991 55526 10025 55538
rect 10545 55526 10579 55538
rect 11099 55526 11133 55538
rect 11653 55526 11687 55538
rect 12207 55526 12241 55538
rect 12761 55526 12795 55538
rect 2211 53550 2212 53574
rect 2292 53550 2293 53574
rect 2765 53550 2766 53574
rect 2846 53550 2847 53574
rect 3319 53550 3320 53574
rect 3400 53550 3401 53574
rect 3873 53550 3874 53574
rect 3954 53550 3955 53574
rect 4427 53550 4428 53574
rect 4508 53550 4509 53574
rect 4981 53550 4982 53574
rect 5062 53550 5063 53574
rect 5535 53550 5536 53574
rect 5616 53550 5617 53574
rect 6089 53550 6090 53574
rect 6170 53550 6171 53574
rect 6643 53550 6644 53574
rect 6724 53550 6725 53574
rect 7197 53550 7198 53574
rect 7278 53550 7279 53574
rect 7751 53550 7752 53574
rect 7832 53550 7833 53574
rect 8305 53550 8306 53574
rect 8386 53550 8387 53574
rect 8859 53550 8860 53574
rect 8940 53550 8941 53574
rect 9413 53550 9414 53574
rect 9494 53550 9495 53574
rect 9967 53550 9968 53574
rect 10048 53550 10049 53574
rect 10521 53550 10522 53574
rect 10602 53550 10603 53574
rect 11075 53550 11076 53574
rect 11156 53550 11157 53574
rect 11629 53550 11630 53574
rect 11710 53550 11711 53574
rect 12183 53550 12184 53574
rect 12264 53550 12265 53574
rect 12737 53550 12738 53574
rect 12818 53550 12819 53574
rect 2235 53526 2269 53538
rect 2789 53526 2823 53538
rect 3343 53526 3377 53538
rect 3897 53526 3931 53538
rect 4451 53526 4485 53538
rect 5005 53526 5039 53538
rect 5559 53526 5593 53538
rect 6113 53526 6147 53538
rect 6667 53526 6701 53538
rect 7221 53526 7255 53538
rect 7775 53526 7809 53538
rect 8329 53526 8363 53538
rect 8883 53526 8917 53538
rect 9437 53526 9471 53538
rect 9991 53526 10025 53538
rect 10545 53526 10579 53538
rect 11099 53526 11133 53538
rect 11653 53526 11687 53538
rect 12207 53526 12241 53538
rect 12761 53526 12795 53538
rect 19352 52294 19402 53694
rect 19502 52294 19630 53694
rect 19658 52294 19786 53694
rect 19814 52294 19942 53694
rect 19970 52294 20098 53694
rect 20126 52294 20254 53694
rect 20282 52294 20410 53694
rect 20438 52294 20566 53694
rect 20594 52294 20722 53694
rect 20750 52294 20878 53694
rect 20906 52294 21034 53694
rect 21062 52294 21190 53694
rect 21218 52294 21346 53694
rect 21374 52294 21502 53694
rect 21530 52294 21658 53694
rect 21686 52294 21814 53694
rect 21842 52294 21970 53694
rect 21998 52294 22126 53694
rect 22154 52294 22282 53694
rect 22310 52294 22438 53694
rect 22466 52294 22594 53694
rect 22622 52294 22750 53694
rect 22778 52294 22906 53694
rect 22934 52294 23062 53694
rect 23090 52294 23218 53694
rect 23246 52294 23374 53694
rect 23402 52294 23530 53694
rect 23558 52294 23686 53694
rect 23714 52294 23842 53694
rect 23870 52294 23998 53694
rect 24026 52294 24154 53694
rect 24182 52294 24310 53694
rect 24338 52294 24466 53694
rect 24494 52294 24622 53694
rect 24650 52294 24778 53694
rect 24806 52294 24934 53694
rect 24962 52294 25090 53694
rect 25118 52294 25246 53694
rect 25274 52294 25402 53694
rect 25430 52294 25558 53694
rect 25586 52294 25714 53694
rect 25742 52294 25870 53694
rect 25898 52294 26026 53694
rect 26054 52294 26182 53694
rect 26210 52294 26338 53694
rect 26366 52294 26494 53694
rect 26522 52294 26650 53694
rect 26678 52294 26806 53694
rect 26834 52294 26962 53694
rect 26990 52294 27118 53694
rect 27146 52294 27196 53694
rect 29067 52850 29117 54250
rect 29217 52850 29345 54250
rect 29373 52850 29501 54250
rect 29529 52850 29657 54250
rect 29685 52850 29813 54250
rect 29841 52850 29969 54250
rect 29997 52850 30125 54250
rect 30153 52850 30281 54250
rect 30309 52850 30437 54250
rect 30465 52850 30593 54250
rect 30621 52850 30749 54250
rect 30777 52850 30905 54250
rect 30933 52850 31061 54250
rect 31089 52850 31217 54250
rect 31245 52850 31373 54250
rect 31401 52850 31451 54250
rect 39130 52488 39180 53888
rect 39280 52488 39408 53888
rect 39436 52488 39564 53888
rect 39592 52488 39720 53888
rect 39748 52488 39876 53888
rect 39904 52488 40032 53888
rect 40060 52488 40188 53888
rect 40216 52488 40344 53888
rect 40372 52488 40500 53888
rect 40528 52488 40656 53888
rect 40684 52488 40812 53888
rect 40840 52488 40968 53888
rect 40996 52488 41124 53888
rect 41152 52488 41280 53888
rect 41308 52488 41436 53888
rect 41464 52488 41592 53888
rect 41620 52488 41748 53888
rect 41776 52488 41904 53888
rect 41932 52488 42060 53888
rect 42088 52488 42216 53888
rect 42244 52488 42372 53888
rect 42400 52488 42528 53888
rect 42556 52488 42684 53888
rect 42712 52488 42840 53888
rect 42868 52488 42996 53888
rect 43024 52488 43152 53888
rect 43180 52488 43308 53888
rect 43336 52488 43464 53888
rect 43492 52488 43620 53888
rect 43648 52488 43776 53888
rect 43804 52488 43932 53888
rect 43960 52488 44088 53888
rect 44116 52488 44244 53888
rect 44272 52488 44400 53888
rect 44428 52488 44556 53888
rect 44584 52488 44712 53888
rect 44740 52488 44868 53888
rect 44896 52488 45024 53888
rect 45052 52488 45180 53888
rect 45208 52488 45336 53888
rect 45364 52488 45492 53888
rect 45520 52488 45648 53888
rect 45676 52488 45804 53888
rect 45832 52488 45960 53888
rect 45988 52488 46116 53888
rect 46144 52488 46272 53888
rect 46300 52488 46428 53888
rect 46456 52488 46584 53888
rect 46612 52488 46740 53888
rect 46768 52488 46896 53888
rect 46924 52488 46974 53888
rect 48845 53044 48895 54444
rect 48995 53044 49123 54444
rect 49151 53044 49279 54444
rect 49307 53044 49435 54444
rect 49463 53044 49591 54444
rect 49619 53044 49747 54444
rect 49775 53044 49903 54444
rect 49931 53044 50059 54444
rect 50087 53044 50215 54444
rect 50243 53044 50371 54444
rect 50399 53044 50527 54444
rect 50555 53044 50683 54444
rect 50711 53044 50839 54444
rect 50867 53044 50995 54444
rect 51023 53044 51151 54444
rect 51179 53044 51229 54444
rect 103638 53996 103710 57996
rect 103909 54029 104027 57963
rect 104298 53996 104358 57996
rect 104558 53996 104630 57996
rect 104829 54029 104947 57963
rect 105218 53996 105278 57996
rect 105478 53996 105550 57996
rect 105749 54029 105867 57963
rect 106138 53996 106198 57996
rect 106398 53996 106470 57996
rect 106669 54029 106787 57963
rect 107058 53996 107118 57996
rect 107318 53996 107390 57996
rect 107589 54029 107707 57963
rect 107978 53996 108038 57996
rect 108238 53996 108310 57996
rect 108509 54029 108627 57963
rect 108898 53996 108958 57996
rect 109158 53996 109230 57996
rect 109429 54029 109547 57963
rect 109818 53996 109878 57996
rect 110078 53996 110150 57996
rect 110349 54029 110467 57963
rect 110738 53996 110798 57996
rect 110998 53996 111070 57996
rect 111269 54029 111387 57963
rect 111658 53996 111718 57996
rect 111918 53996 111990 57996
rect 112189 54029 112307 57963
rect 112578 53996 112638 57996
rect 112838 53996 112910 57996
rect 113109 54029 113227 57963
rect 113498 53996 113558 57996
rect 127615 55792 127617 55917
rect 62707 53804 62708 53828
rect 62788 53804 62789 53828
rect 63261 53804 63262 53828
rect 63342 53804 63343 53828
rect 63815 53804 63816 53828
rect 63896 53804 63897 53828
rect 64369 53804 64370 53828
rect 64450 53804 64451 53828
rect 64923 53804 64924 53828
rect 65004 53804 65005 53828
rect 65477 53804 65478 53828
rect 65558 53804 65559 53828
rect 66031 53804 66032 53828
rect 66112 53804 66113 53828
rect 66585 53804 66586 53828
rect 66666 53804 66667 53828
rect 67139 53804 67140 53828
rect 67220 53804 67221 53828
rect 67693 53804 67694 53828
rect 67774 53804 67775 53828
rect 68247 53804 68248 53828
rect 68328 53804 68329 53828
rect 68801 53804 68802 53828
rect 68882 53804 68883 53828
rect 69355 53804 69356 53828
rect 69436 53804 69437 53828
rect 69909 53804 69910 53828
rect 69990 53804 69991 53828
rect 70463 53804 70464 53828
rect 70544 53804 70545 53828
rect 71017 53804 71018 53828
rect 71098 53804 71099 53828
rect 71571 53804 71572 53828
rect 71652 53804 71653 53828
rect 72125 53804 72126 53828
rect 72206 53804 72207 53828
rect 72679 53804 72680 53828
rect 72760 53804 72761 53828
rect 73233 53804 73234 53828
rect 73314 53804 73315 53828
rect 62731 53780 62765 53792
rect 63285 53780 63319 53792
rect 63839 53780 63873 53792
rect 64393 53780 64427 53792
rect 64947 53780 64981 53792
rect 65501 53780 65535 53792
rect 66055 53780 66089 53792
rect 66609 53780 66643 53792
rect 67163 53780 67197 53792
rect 67717 53780 67751 53792
rect 68271 53780 68305 53792
rect 68825 53780 68859 53792
rect 69379 53780 69413 53792
rect 69933 53780 69967 53792
rect 70487 53780 70521 53792
rect 71041 53780 71075 53792
rect 71595 53780 71629 53792
rect 72149 53780 72183 53792
rect 72703 53780 72737 53792
rect 73257 53780 73291 53792
rect 81709 53610 81710 53634
rect 81790 53610 81791 53634
rect 82263 53610 82264 53634
rect 82344 53610 82345 53634
rect 82817 53610 82818 53634
rect 82898 53610 82899 53634
rect 83371 53610 83372 53634
rect 83452 53610 83453 53634
rect 83925 53610 83926 53634
rect 84006 53610 84007 53634
rect 84479 53610 84480 53634
rect 84560 53610 84561 53634
rect 85033 53610 85034 53634
rect 85114 53610 85115 53634
rect 85587 53610 85588 53634
rect 85668 53610 85669 53634
rect 86141 53610 86142 53634
rect 86222 53610 86223 53634
rect 86695 53610 86696 53634
rect 86776 53610 86777 53634
rect 87249 53610 87250 53634
rect 87330 53610 87331 53634
rect 87803 53610 87804 53634
rect 87884 53610 87885 53634
rect 88357 53610 88358 53634
rect 88438 53610 88439 53634
rect 88911 53610 88912 53634
rect 88992 53610 88993 53634
rect 89465 53610 89466 53634
rect 89546 53610 89547 53634
rect 90019 53610 90020 53634
rect 90100 53610 90101 53634
rect 90573 53610 90574 53634
rect 90654 53610 90655 53634
rect 91127 53610 91128 53634
rect 91208 53610 91209 53634
rect 91681 53610 91682 53634
rect 91762 53610 91763 53634
rect 92235 53610 92236 53634
rect 92316 53610 92317 53634
rect 81733 53586 81767 53598
rect 82287 53586 82321 53598
rect 82841 53586 82875 53598
rect 83395 53586 83429 53598
rect 83949 53586 83983 53598
rect 84503 53586 84537 53598
rect 85057 53586 85091 53598
rect 85611 53586 85645 53598
rect 86165 53586 86199 53598
rect 86719 53586 86753 53598
rect 87273 53586 87307 53598
rect 87827 53586 87861 53598
rect 88381 53586 88415 53598
rect 88935 53586 88969 53598
rect 89489 53586 89523 53598
rect 90043 53586 90077 53598
rect 90597 53586 90631 53598
rect 91151 53586 91185 53598
rect 91705 53586 91739 53598
rect 92259 53586 92293 53598
rect 2211 51550 2212 51574
rect 2292 51550 2293 51574
rect 2765 51550 2766 51574
rect 2846 51550 2847 51574
rect 3319 51550 3320 51574
rect 3400 51550 3401 51574
rect 3873 51550 3874 51574
rect 3954 51550 3955 51574
rect 4427 51550 4428 51574
rect 4508 51550 4509 51574
rect 4981 51550 4982 51574
rect 5062 51550 5063 51574
rect 5535 51550 5536 51574
rect 5616 51550 5617 51574
rect 6089 51550 6090 51574
rect 6170 51550 6171 51574
rect 6643 51550 6644 51574
rect 6724 51550 6725 51574
rect 7197 51550 7198 51574
rect 7278 51550 7279 51574
rect 7751 51550 7752 51574
rect 7832 51550 7833 51574
rect 8305 51550 8306 51574
rect 8386 51550 8387 51574
rect 8859 51550 8860 51574
rect 8940 51550 8941 51574
rect 9413 51550 9414 51574
rect 9494 51550 9495 51574
rect 9967 51550 9968 51574
rect 10048 51550 10049 51574
rect 10521 51550 10522 51574
rect 10602 51550 10603 51574
rect 11075 51550 11076 51574
rect 11156 51550 11157 51574
rect 11629 51550 11630 51574
rect 11710 51550 11711 51574
rect 12183 51550 12184 51574
rect 12264 51550 12265 51574
rect 12737 51550 12738 51574
rect 12818 51550 12819 51574
rect 2235 51526 2269 51538
rect 2789 51526 2823 51538
rect 3343 51526 3377 51538
rect 3897 51526 3931 51538
rect 4451 51526 4485 51538
rect 5005 51526 5039 51538
rect 5559 51526 5593 51538
rect 6113 51526 6147 51538
rect 6667 51526 6701 51538
rect 7221 51526 7255 51538
rect 7775 51526 7809 51538
rect 8329 51526 8363 51538
rect 8883 51526 8917 51538
rect 9437 51526 9471 51538
rect 9991 51526 10025 51538
rect 10545 51526 10579 51538
rect 11099 51526 11133 51538
rect 11653 51526 11687 51538
rect 12207 51526 12241 51538
rect 12761 51526 12795 51538
rect 29647 50763 29697 51763
rect 30497 50763 30547 51763
rect 30799 50763 30849 51763
rect 31649 50763 31699 51763
rect 49425 50957 49475 51957
rect 50275 50957 50325 51957
rect 50577 50957 50627 51957
rect 51427 50957 51477 51957
rect 62707 51804 62708 51828
rect 62788 51804 62789 51828
rect 63261 51804 63262 51828
rect 63342 51804 63343 51828
rect 63815 51804 63816 51828
rect 63896 51804 63897 51828
rect 64369 51804 64370 51828
rect 64450 51804 64451 51828
rect 64923 51804 64924 51828
rect 65004 51804 65005 51828
rect 65477 51804 65478 51828
rect 65558 51804 65559 51828
rect 66031 51804 66032 51828
rect 66112 51804 66113 51828
rect 66585 51804 66586 51828
rect 66666 51804 66667 51828
rect 67139 51804 67140 51828
rect 67220 51804 67221 51828
rect 67693 51804 67694 51828
rect 67774 51804 67775 51828
rect 68247 51804 68248 51828
rect 68328 51804 68329 51828
rect 68801 51804 68802 51828
rect 68882 51804 68883 51828
rect 69355 51804 69356 51828
rect 69436 51804 69437 51828
rect 69909 51804 69910 51828
rect 69990 51804 69991 51828
rect 70463 51804 70464 51828
rect 70544 51804 70545 51828
rect 71017 51804 71018 51828
rect 71098 51804 71099 51828
rect 71571 51804 71572 51828
rect 71652 51804 71653 51828
rect 72125 51804 72126 51828
rect 72206 51804 72207 51828
rect 72679 51804 72680 51828
rect 72760 51804 72761 51828
rect 73233 51804 73234 51828
rect 73314 51804 73315 51828
rect 62731 51780 62765 51792
rect 63285 51780 63319 51792
rect 63839 51780 63873 51792
rect 64393 51780 64427 51792
rect 64947 51780 64981 51792
rect 65501 51780 65535 51792
rect 66055 51780 66089 51792
rect 66609 51780 66643 51792
rect 67163 51780 67197 51792
rect 67717 51780 67751 51792
rect 68271 51780 68305 51792
rect 68825 51780 68859 51792
rect 69379 51780 69413 51792
rect 69933 51780 69967 51792
rect 70487 51780 70521 51792
rect 71041 51780 71075 51792
rect 71595 51780 71629 51792
rect 72149 51780 72183 51792
rect 72703 51780 72737 51792
rect 73257 51780 73291 51792
rect 81709 51610 81710 51634
rect 81790 51610 81791 51634
rect 82263 51610 82264 51634
rect 82344 51610 82345 51634
rect 82817 51610 82818 51634
rect 82898 51610 82899 51634
rect 83371 51610 83372 51634
rect 83452 51610 83453 51634
rect 83925 51610 83926 51634
rect 84006 51610 84007 51634
rect 84479 51610 84480 51634
rect 84560 51610 84561 51634
rect 85033 51610 85034 51634
rect 85114 51610 85115 51634
rect 85587 51610 85588 51634
rect 85668 51610 85669 51634
rect 86141 51610 86142 51634
rect 86222 51610 86223 51634
rect 86695 51610 86696 51634
rect 86776 51610 86777 51634
rect 87249 51610 87250 51634
rect 87330 51610 87331 51634
rect 87803 51610 87804 51634
rect 87884 51610 87885 51634
rect 88357 51610 88358 51634
rect 88438 51610 88439 51634
rect 88911 51610 88912 51634
rect 88992 51610 88993 51634
rect 89465 51610 89466 51634
rect 89546 51610 89547 51634
rect 90019 51610 90020 51634
rect 90100 51610 90101 51634
rect 90573 51610 90574 51634
rect 90654 51610 90655 51634
rect 91127 51610 91128 51634
rect 91208 51610 91209 51634
rect 91681 51610 91682 51634
rect 91762 51610 91763 51634
rect 92235 51610 92236 51634
rect 92316 51610 92317 51634
rect 81733 51586 81767 51598
rect 82287 51586 82321 51598
rect 82841 51586 82875 51598
rect 83395 51586 83429 51598
rect 83949 51586 83983 51598
rect 84503 51586 84537 51598
rect 85057 51586 85091 51598
rect 85611 51586 85645 51598
rect 86165 51586 86199 51598
rect 86719 51586 86753 51598
rect 87273 51586 87307 51598
rect 87827 51586 87861 51598
rect 88381 51586 88415 51598
rect 88935 51586 88969 51598
rect 89489 51586 89523 51598
rect 90043 51586 90077 51598
rect 90597 51586 90631 51598
rect 91151 51586 91185 51598
rect 91705 51586 91739 51598
rect 92259 51586 92293 51598
rect -432 50006 -366 50022
rect 6799 49836 6885 49872
rect 3431 49642 3783 49668
rect 4255 49642 4607 49668
rect 5079 49642 5431 49668
rect 5903 49642 6255 49668
rect 3457 46643 3458 49642
rect 3757 46643 3783 49642
rect 3457 46642 3783 46643
rect 4281 46643 4282 49642
rect 4581 46643 4607 49642
rect 4281 46642 4607 46643
rect 5105 46643 5106 49642
rect 5405 46643 5431 49642
rect 5105 46642 5431 46643
rect 5929 46643 5930 49642
rect 6229 46643 6255 49642
rect 5929 46642 6255 46643
rect 6799 46448 6835 49836
rect 6849 46448 6885 49836
rect 7429 49642 7781 49668
rect 8253 49642 8605 49668
rect 9077 49642 9429 49668
rect 9901 49642 10253 49668
rect 7455 46643 7456 49642
rect 7755 46643 7781 49642
rect 7455 46642 7781 46643
rect 8279 46643 8280 49642
rect 8579 46643 8605 49642
rect 8279 46642 8605 46643
rect 9103 46643 9104 49642
rect 9403 46643 9429 49642
rect 9103 46642 9429 46643
rect 9927 46643 9928 49642
rect 10227 46643 10253 49642
rect 21039 49519 21089 50519
rect 21889 49519 21939 50519
rect 22191 49519 22241 50519
rect 23841 49519 23891 50519
rect 24143 49519 24193 50519
rect 25793 49519 25843 50519
rect 26095 49519 26145 50519
rect 27745 49519 27795 50519
rect 28047 49519 28097 50519
rect 29697 49519 29747 50519
rect 29999 49519 30049 50519
rect 31649 49519 31699 50519
rect 40817 49713 40867 50713
rect 41667 49713 41717 50713
rect 41969 49713 42019 50713
rect 43619 49713 43669 50713
rect 43921 49713 43971 50713
rect 45571 49713 45621 50713
rect 45873 49713 45923 50713
rect 47523 49713 47573 50713
rect 47825 49713 47875 50713
rect 49475 49713 49525 50713
rect 49777 49713 49827 50713
rect 51427 49713 51477 50713
rect 101758 50520 101808 51920
rect 101908 50520 102036 51920
rect 102064 50520 102192 51920
rect 102220 50520 102348 51920
rect 102376 50520 102504 51920
rect 102532 50520 102660 51920
rect 102688 50520 102816 51920
rect 102844 50520 102972 51920
rect 103000 50520 103128 51920
rect 103156 50520 103284 51920
rect 103312 50520 103440 51920
rect 103468 50520 103596 51920
rect 103624 50520 103752 51920
rect 103780 50520 103908 51920
rect 103936 50520 104064 51920
rect 104092 50520 104220 51920
rect 104248 50520 104376 51920
rect 104404 50520 104532 51920
rect 104560 50520 104688 51920
rect 104716 50520 104844 51920
rect 104872 50520 105000 51920
rect 105028 50520 105156 51920
rect 105184 50520 105312 51920
rect 105340 50520 105468 51920
rect 105496 50520 105624 51920
rect 105652 50520 105780 51920
rect 105808 50520 105936 51920
rect 105964 50520 106092 51920
rect 106120 50520 106248 51920
rect 106276 50520 106404 51920
rect 106432 50520 106560 51920
rect 106588 50520 106716 51920
rect 106744 50520 106872 51920
rect 106900 50520 107028 51920
rect 107056 50520 107184 51920
rect 107212 50520 107340 51920
rect 107368 50520 107496 51920
rect 107524 50520 107652 51920
rect 107680 50520 107808 51920
rect 107836 50520 107964 51920
rect 107992 50520 108120 51920
rect 108148 50520 108276 51920
rect 108304 50520 108432 51920
rect 108460 50520 108588 51920
rect 108616 50520 108744 51920
rect 108772 50520 108900 51920
rect 108928 50520 109056 51920
rect 109084 50520 109212 51920
rect 109240 50520 109368 51920
rect 109396 50520 109524 51920
rect 109552 50520 109602 51920
rect 111473 51076 111523 52476
rect 111623 51076 111751 52476
rect 111779 51076 111907 52476
rect 111935 51076 112063 52476
rect 112091 51076 112219 52476
rect 112247 51076 112375 52476
rect 112403 51076 112531 52476
rect 112559 51076 112687 52476
rect 112715 51076 112843 52476
rect 112871 51076 112999 52476
rect 113027 51076 113155 52476
rect 113183 51076 113311 52476
rect 113339 51076 113467 52476
rect 113495 51076 113623 52476
rect 113651 51076 113779 52476
rect 113807 51076 113857 52476
rect 62707 49804 62708 49828
rect 62788 49804 62789 49828
rect 63261 49804 63262 49828
rect 63342 49804 63343 49828
rect 63815 49804 63816 49828
rect 63896 49804 63897 49828
rect 64369 49804 64370 49828
rect 64450 49804 64451 49828
rect 64923 49804 64924 49828
rect 65004 49804 65005 49828
rect 65477 49804 65478 49828
rect 65558 49804 65559 49828
rect 66031 49804 66032 49828
rect 66112 49804 66113 49828
rect 66585 49804 66586 49828
rect 66666 49804 66667 49828
rect 67139 49804 67140 49828
rect 67220 49804 67221 49828
rect 67693 49804 67694 49828
rect 67774 49804 67775 49828
rect 68247 49804 68248 49828
rect 68328 49804 68329 49828
rect 68801 49804 68802 49828
rect 68882 49804 68883 49828
rect 69355 49804 69356 49828
rect 69436 49804 69437 49828
rect 69909 49804 69910 49828
rect 69990 49804 69991 49828
rect 70463 49804 70464 49828
rect 70544 49804 70545 49828
rect 71017 49804 71018 49828
rect 71098 49804 71099 49828
rect 71571 49804 71572 49828
rect 71652 49804 71653 49828
rect 72125 49804 72126 49828
rect 72206 49804 72207 49828
rect 72679 49804 72680 49828
rect 72760 49804 72761 49828
rect 73233 49804 73234 49828
rect 73314 49804 73315 49828
rect 62731 49780 62765 49792
rect 63285 49780 63319 49792
rect 63839 49780 63873 49792
rect 64393 49780 64427 49792
rect 64947 49780 64981 49792
rect 65501 49780 65535 49792
rect 66055 49780 66089 49792
rect 66609 49780 66643 49792
rect 67163 49780 67197 49792
rect 67717 49780 67751 49792
rect 68271 49780 68305 49792
rect 68825 49780 68859 49792
rect 69379 49780 69413 49792
rect 69933 49780 69967 49792
rect 70487 49780 70521 49792
rect 71041 49780 71075 49792
rect 71595 49780 71629 49792
rect 72149 49780 72183 49792
rect 72703 49780 72737 49792
rect 73257 49780 73291 49792
rect 81709 49610 81710 49634
rect 81790 49610 81791 49634
rect 82263 49610 82264 49634
rect 82344 49610 82345 49634
rect 82817 49610 82818 49634
rect 82898 49610 82899 49634
rect 83371 49610 83372 49634
rect 83452 49610 83453 49634
rect 83925 49610 83926 49634
rect 84006 49610 84007 49634
rect 84479 49610 84480 49634
rect 84560 49610 84561 49634
rect 85033 49610 85034 49634
rect 85114 49610 85115 49634
rect 85587 49610 85588 49634
rect 85668 49610 85669 49634
rect 86141 49610 86142 49634
rect 86222 49610 86223 49634
rect 86695 49610 86696 49634
rect 86776 49610 86777 49634
rect 87249 49610 87250 49634
rect 87330 49610 87331 49634
rect 87803 49610 87804 49634
rect 87884 49610 87885 49634
rect 88357 49610 88358 49634
rect 88438 49610 88439 49634
rect 88911 49610 88912 49634
rect 88992 49610 88993 49634
rect 89465 49610 89466 49634
rect 89546 49610 89547 49634
rect 90019 49610 90020 49634
rect 90100 49610 90101 49634
rect 90573 49610 90574 49634
rect 90654 49610 90655 49634
rect 91127 49610 91128 49634
rect 91208 49610 91209 49634
rect 91681 49610 91682 49634
rect 91762 49610 91763 49634
rect 92235 49610 92236 49634
rect 92316 49610 92317 49634
rect 81733 49586 81767 49598
rect 82287 49586 82321 49598
rect 82841 49586 82875 49598
rect 83395 49586 83429 49598
rect 83949 49586 83983 49598
rect 84503 49586 84537 49598
rect 85057 49586 85091 49598
rect 85611 49586 85645 49598
rect 86165 49586 86199 49598
rect 86719 49586 86753 49598
rect 87273 49586 87307 49598
rect 87827 49586 87861 49598
rect 88381 49586 88415 49598
rect 88935 49586 88969 49598
rect 89489 49586 89523 49598
rect 90043 49586 90077 49598
rect 90597 49586 90631 49598
rect 91151 49586 91185 49598
rect 91705 49586 91739 49598
rect 92259 49586 92293 49598
rect 21039 48275 21089 49275
rect 21889 48275 21939 49275
rect 22191 48275 22241 49275
rect 23841 48275 23891 49275
rect 24143 48275 24193 49275
rect 25793 48275 25843 49275
rect 26095 48275 26145 49275
rect 27745 48275 27795 49275
rect 28047 48275 28097 49275
rect 29697 48275 29747 49275
rect 29999 48275 30049 49275
rect 31649 48275 31699 49275
rect 40817 48469 40867 49469
rect 41667 48469 41717 49469
rect 41969 48469 42019 49469
rect 43619 48469 43669 49469
rect 43921 48469 43971 49469
rect 45571 48469 45621 49469
rect 45873 48469 45923 49469
rect 47523 48469 47573 49469
rect 47825 48469 47875 49469
rect 49475 48469 49525 49469
rect 49777 48469 49827 49469
rect 51427 48469 51477 49469
rect 112053 48989 112103 49989
rect 112903 48989 112953 49989
rect 113205 48989 113255 49989
rect 114055 48989 114105 49989
rect 60064 48260 60130 48276
rect 21039 47031 21089 48031
rect 21889 47031 21939 48031
rect 22191 47031 22241 48031
rect 23841 47031 23891 48031
rect 24143 47031 24193 48031
rect 25793 47031 25843 48031
rect 26095 47031 26145 48031
rect 27745 47031 27795 48031
rect 28047 47031 28097 48031
rect 29697 47031 29747 48031
rect 29999 47031 30049 48031
rect 31649 47031 31699 48031
rect 40817 47225 40867 48225
rect 41667 47225 41717 48225
rect 41969 47225 42019 48225
rect 43619 47225 43669 48225
rect 43921 47225 43971 48225
rect 45571 47225 45621 48225
rect 45873 47225 45923 48225
rect 47523 47225 47573 48225
rect 47825 47225 47875 48225
rect 49475 47225 49525 48225
rect 49777 47225 49827 48225
rect 51427 47225 51477 48225
rect 67295 48090 67381 48126
rect 63927 47896 64279 47922
rect 64751 47896 65103 47922
rect 65575 47896 65927 47922
rect 66399 47896 66751 47922
rect 9927 46642 10253 46643
rect 6799 46412 6885 46448
rect 63953 44897 63954 47896
rect 64253 44897 64279 47896
rect 63953 44896 64279 44897
rect 64777 44897 64778 47896
rect 65077 44897 65103 47896
rect 64777 44896 65103 44897
rect 65601 44897 65602 47896
rect 65901 44897 65927 47896
rect 65601 44896 65927 44897
rect 66425 44897 66426 47896
rect 66725 44897 66751 47896
rect 66425 44896 66751 44897
rect 67295 44702 67331 48090
rect 67345 44702 67381 48090
rect 79066 48066 79132 48082
rect 67925 47896 68277 47922
rect 68749 47896 69101 47922
rect 69573 47896 69925 47922
rect 70397 47896 70749 47922
rect 67951 44897 67952 47896
rect 68251 44897 68277 47896
rect 67951 44896 68277 44897
rect 68775 44897 68776 47896
rect 69075 44897 69101 47896
rect 68775 44896 69101 44897
rect 69599 44897 69600 47896
rect 69899 44897 69925 47896
rect 69599 44896 69925 44897
rect 70423 44897 70424 47896
rect 70723 44897 70749 47896
rect 86297 47896 86383 47932
rect 82929 47702 83281 47728
rect 83753 47702 84105 47728
rect 84577 47702 84929 47728
rect 85401 47702 85753 47728
rect 70423 44896 70749 44897
rect 82955 44703 82956 47702
rect 83255 44703 83281 47702
rect 82955 44702 83281 44703
rect 83779 44703 83780 47702
rect 84079 44703 84105 47702
rect 83779 44702 84105 44703
rect 84603 44703 84604 47702
rect 84903 44703 84929 47702
rect 84603 44702 84929 44703
rect 85427 44703 85428 47702
rect 85727 44703 85753 47702
rect 85427 44702 85753 44703
rect 67295 44666 67381 44702
rect 86297 44508 86333 47896
rect 86347 44508 86383 47896
rect 103445 47745 103495 48745
rect 104295 47745 104345 48745
rect 104597 47745 104647 48745
rect 106247 47745 106297 48745
rect 106549 47745 106599 48745
rect 108199 47745 108249 48745
rect 108501 47745 108551 48745
rect 110151 47745 110201 48745
rect 110453 47745 110503 48745
rect 112103 47745 112153 48745
rect 112405 47745 112455 48745
rect 114055 47745 114105 48745
rect 86927 47702 87279 47728
rect 87751 47702 88103 47728
rect 88575 47702 88927 47728
rect 89399 47702 89751 47728
rect 86953 44703 86954 47702
rect 87253 44703 87279 47702
rect 86953 44702 87279 44703
rect 87777 44703 87778 47702
rect 88077 44703 88103 47702
rect 87777 44702 88103 44703
rect 88601 44703 88602 47702
rect 88901 44703 88927 47702
rect 88601 44702 88927 44703
rect 89425 44703 89426 47702
rect 89725 44703 89751 47702
rect 103445 46501 103495 47501
rect 104295 46501 104345 47501
rect 104597 46501 104647 47501
rect 106247 46501 106297 47501
rect 106549 46501 106599 47501
rect 108199 46501 108249 47501
rect 108501 46501 108551 47501
rect 110151 46501 110201 47501
rect 110453 46501 110503 47501
rect 112103 46501 112153 47501
rect 112405 46501 112455 47501
rect 114055 46501 114105 47501
rect 103445 45257 103495 46257
rect 104295 45257 104345 46257
rect 104597 45257 104647 46257
rect 106247 45257 106297 46257
rect 106549 45257 106599 46257
rect 108199 45257 108249 46257
rect 108501 45257 108551 46257
rect 110151 45257 110201 46257
rect 110453 45257 110503 46257
rect 112103 45257 112153 46257
rect 112405 45257 112455 46257
rect 114055 45257 114105 46257
rect 89425 44702 89751 44703
rect 86297 44472 86383 44508
use sky130_ef_io__vdda_lvc_pad  sky130_ef_io__vdda_lvc_pad_0
timestamp 1584383356
transform 1 0 -868 0 1 91931
box 0 -61 15000 39593
use sky130_ef_io__vdda_hvc_pad  sky130_ef_io__vdda_hvc_pad_0
timestamp 1584383356
transform 1 0 19686 0 1 92471
box 0 -407 15000 39593
use sky130_ef_io__vccd_lvc_pad  sky130_ef_io__vccd_lvc_pad_0
timestamp 1584383356
transform 1 0 38106 0 1 91155
box 0 -61 15000 39593
use sky130_ef_io__vccd_hvc_pad  sky130_ef_io__vccd_hvc_pad_0
timestamp 1584383356
transform 1 0 56526 0 1 91335
box 0 -435 15000 39593
use sky130_ef_io__vddio_hvc_pad  sky130_ef_io__vddio_hvc_pad_0
timestamp 1584383356
transform 1 0 77078 0 1 92305
box 0 -435 15000 39593
use sky130_ef_io__vddio_lvc_pad  sky130_ef_io__vddio_lvc_pad_0
timestamp 1584383356
transform 1 0 97048 0 1 92319
box 0 -61 15000 39593
use sky130_ef_io__gpiov2_pad  sky130_ef_io__gpiov2_pad_0
timestamp 1584383356
transform 1 0 119295 0 1 92724
box -143 -466 16134 39593
use sky130_ef_io__top_xres4v2  sky130_ef_io__top_xres4v2_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1584046481
transform 1 0 140197 0 1 92452
box -103 0 15124 40000
use sky130_ef_io__top_gpio_ovtv2  sky130_ef_io__top_gpio_ovtv2_0 ~/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_io/mag
timestamp 1584046481
transform 1 0 160920 0 1 92540
box -80 -88 28211 40076
use sky130_ef_io__vssd_lvc_pad  sky130_ef_io__vssd_lvc_pad_0
timestamp 1584383356
transform 1 0 -480 0 1 46173
box 0 -61 15000 39593
use sky130_ef_io__vssd_hvc_pad  sky130_ef_io__vssd_hvc_pad_0
timestamp 1584383356
transform 1 0 18134 0 1 46741
box 0 -435 15000 39593
use sky130_ef_io__vssa_hvc_pad  sky130_ef_io__vssa_hvc_pad_0
timestamp 1584383356
transform 1 0 37912 0 1 46935
box 0 -435 15000 39593
use sky130_ef_io__vssa_lvc_pad  sky130_ef_io__vssa_lvc_pad_0
timestamp 1584383356
transform 1 0 60016 0 1 44427
box 0 -61 15000 39593
use sky130_ef_io__vssio_lvc_pad  sky130_ef_io__vssio_lvc_pad_0
timestamp 1584383356
transform 1 0 79018 0 1 44233
box 0 -61 15000 39593
use sky130_ef_io__vssio_hvc_pad  sky130_ef_io__vssio_hvc_pad_0
timestamp 1584383356
transform 1 0 100540 0 1 44967
box 0 -407 15000 39593
use sky130_ef_io__corner_pad  sky130_ef_io__corner_pad_0
timestamp 1584383356
transform 1 0 123795 0 1 46420
box -181 -114 40000 40800
<< end >>
